module physics_coprocessor(
	clock, reset, 			// Master clock, reset signals

	mass_in, gravity_in, wind_in, 	// Constants set for the player
	start_Position, 		// Starting position [x, y]

	controller_in, 			// Input from controller joystick
	knockback_in,			// Input from attack coprocessor
	attack_in,				// Input from attack coprocessor


	wall, 					// Hitting walls

	freeze_in,				// Holds player still

	position 				// Output position [x, y]
);

	// Inputs
	input clock, reset;
	input [31:0] mass_in, gravity_in, wind_in;
	input [31:0] start_Position;
	input [31:0] controller_in, knockback_in;
	input [31:0] wall;
	input attack_in;
	input freeze_in;

	// Output Position
	output [31:0] position;

	// Input from Controller
	wire signed [8:0] joystick_x, joystick_y; // Unsigned values from 0 to 255 representing joystick position
	assign joystick_x[7:0] = controller_in[15:8];
	assign joystick_x[8] = 1'b0;
	assign joystick_y[7:0] = controller_in[7:0];
	assign joystick_y[8] = 1'b0;
	wire jump;
	wire platform_Thru;
	assign jump = joystick_y[7] & joystick_y[6] & joystick_y[5] & joystick_y[4]; // Joystick Y 240 to 255 (up)
	assign platform_Thru = ~joystick_y[7] & ~joystick_y[6] & ~joystick_y[5] & ~joystick_y[4]; // Joystick Y 0 to 15 (down)
	
	// Input from Collisions
	wire wall_Left, wall_Right, wall_Up, wall_Down, platform_Down;
	assign wall_Left = wall[3];
	assign wall_Right = wall[2];
	assign wall_Up = wall[0];
	assign wall_Down = wall[1];
	assign platform_Down = wall[4];

	// Input Physics Parameters
	wire [47:0] mass, gravity, wind;
	wire signed [47:0] move_x, move_y, knockback_x, knockback_y;
	assign mass[31:0] = mass_in;
	assign mass[47:32] = 16'b0;
	assign gravity[31:0] = gravity_in;
	assign gravity[47:32] = 16'b0;
	assign wind[31:0] = wind_in;
	assign wind[47:32] = 16'b0;
	assign move_x[16:8] = joystick_x - 9'b001110000; // Map joystick values to -128 to 127
	assign move_x[7:0] = 8'b0;
	assign move_y[16:8] = joystick_y - 9'b001110000; // Map joystick values to -128 to 127
	assign move_y[7:0] = 8'b0;
	assign knockback_x[15:0] = knockback_in[31:16]; // Split knockback into x, y
	assign knockback_y[15:0] = knockback_in[15:0];
	genvar i;
	generate // Extend joystick, knockback values to 32 bit signed values
		for(i = 17; i < 48; i = i + 1) begin: signextend1
			assign move_x[i] = move_x[16];
			assign move_y[i] = move_y[16];
		end
		for(i = 16; i < 48; i = i + 1) begin: signextend2
			assign knockback_x[i] = knockback_in[31];
			assign knockback_y[i] = knockback_in[15];
		end
	endgenerate

	 // X, Y position components
    reg [47:0] pos_x, pos_y;

    // Stored Values
    reg signed [47:0] vel_x, vel_y;
    reg signed [47:0] accel_x, accel_y;

    // Vibration Values
    reg [47:0] vibr_pos_y;
    wire vibr_dir;
    assign vibr_dir = (pos_y < vibr_pos_y + 48'd10000000)? 1'b1 : 1'b0;

    // Attack start, end value
    reg attack_prev;

    // Separate input, output components
    assign position[31:16] = pos_x[47:32];
    assign position[15:0] = pos_y[47:32];

    // Update values every cycle
    always@(posedge clock) begin
	 
		// Reset
		if(reset) begin
		   accel_x <= 48'b0;
			accel_y <= 48'b0;
			vel_x <= 48'b0;
			vel_y <= 48'b0;
			pos_x [47:32] <= start_Position[31:16];
			pos_x [31:0] <= 32'b0;
			pos_y [47:32] <= start_Position[15:0];
			pos_y [31:0] <= 32'b0;
		end

    	// Acceleration, velocity update for in air
    	else if(~freeze_in & ~attack_in & ~wall_Down & ~platform_Down) begin
    		accel_x <= move_x / mass;// - vel_x * vel_x * vel_x / wind;
    		accel_y <= move_y / mass - gravity;// - vel_y * vel_y * vel_y / wind;
    		vel_x <= move_x / mass; // TODO Fix for Collisions L, R
    		if(~jump) vel_y <= move_y / mass - gravity; // TODO Fix for collisions U, jumps
			else vel_y <= move_y / mass;
    		pos_x <= pos_x + vel_x;
    		pos_y <= pos_y + vel_y;
    	end

    	// Acceleration, velocity update for on ground
    	else if(~freeze_in & ~attack_in & (wall_Down | platform_Down)) begin
    		accel_x <= 48'b0;
    		accel_y <= 48'b0;
    		vel_x <= move_x / mass; // TODO Fix for Collisions L, R
    		if(~jump) vel_y <= 48'b0; // TODO Fix for platform thru, jumps
			else vel_y <= move_y / mass;
    		pos_x <= pos_x + vel_x;
    	end

    	// Start of attack
    	if(~reset & attack_in & ~attack_prev) begin
    		attack_prev <= attack_in;
	    	vibr_pos_y <= pos_y + 48'h00010000; // Start up 1 pixel to be off the ground
	    	pos_y <= pos_y + 48'h00010000;
	    end

    	// During Attack
    	if(~reset & attack_prev) begin
    		accel_x <= 48'b0;
	    	accel_y <= 48'b0;
	    	attack_prev <= attack_in;
    		// Knockback velocity
    		vel_x <= knockback_x / mass;
	    	vel_y <= knockback_y / mass;
     		// Attack vibration
    		if(vibr_dir)
    			pos_y <= pos_y + 48'd2;
    		else
    			pos_y <= pos_y - 48'd2; 
    	end

    end

endmodule
