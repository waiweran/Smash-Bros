module multiplier(inA, inB, out);
	input [31:0] inA, inB;
	output [63:0] out;

	wire wire129, wire130, wire131, wire132, wire133, wire134, wire135, wire136, wire137, wire138, wire139, wire140, wire141, wire142, wire143, wire144, wire145, wire146, wire147, wire148, wire149, wire150, wire151, wire152, wire153, wire154, wire155, wire156, wire157, wire158, wire159, wire160, wire161, wire162, wire163, wire164, wire165, wire166, wire167, wire168, wire169, wire170, wire171, wire172, wire173, wire174, wire175, wire176, wire177, wire178, wire179, wire180, wire181, wire182, wire183, wire184, wire185, wire186, wire187, wire188, wire189, wire190, wire191, wire192, wire193, wire194, wire195, wire196, wire197, wire198, wire199, wire200, wire201, wire202, wire203, wire204, wire205, wire206, wire207, wire208, wire209, wire210, wire211, wire212, wire213, wire214, wire215, wire216, wire217, wire218, wire219, wire220, wire221, wire222, wire223, wire224, wire225, wire226, wire227, wire228, wire229, wire230, wire231, wire232, wire233, wire234, wire235, wire236, wire237, wire238, wire239, wire240, wire241, wire242, wire243, wire244, wire245, wire246, wire247, wire248, wire249, wire250, wire251, wire252, wire253, wire254, wire255, wire256, wire257, wire258, wire259, wire260, wire261, wire262, wire263, wire264, wire265, wire266, wire267, wire268, wire269, wire270, wire271, wire272, wire273, wire274, wire275, wire276, wire277, wire278, wire279, wire280, wire281, wire282, wire283, wire284, wire285, wire286, wire287, wire288, wire289, wire290, wire291, wire292, wire293, wire294, wire295, wire296, wire297, wire298, wire299, wire300, wire301, wire302, wire303, wire304, wire305, wire306, wire307, wire308, wire309, wire310, wire311, wire312, wire313, wire314, wire315, wire316, wire317, wire318, wire319, wire320, wire321, wire322, wire323, wire324, wire325, wire326, wire327, wire328, wire329, wire330, wire331, wire332, wire333, wire334, wire335, wire336, wire337, wire338, wire339, wire340, wire341, wire342, wire343, wire344, wire345, wire346, wire347, wire348, wire349, wire350, wire351, wire352, wire353, wire354, wire355, wire356, wire357, wire358, wire359, wire360, wire361, wire362, wire363, wire364, wire365, wire366, wire367, wire368, wire369, wire370, wire371, wire372, wire373, wire374, wire375, wire376, wire377, wire378, wire379, wire380, wire381, wire382, wire383, wire384, wire385, wire386, wire387, wire388, wire389, wire390, wire391, wire392, wire393, wire394, wire395, wire396, wire397, wire398, wire399, wire400, wire401, wire402, wire403, wire404, wire405, wire406, wire407, wire408, wire409, wire410, wire411, wire412, wire413, wire414, wire415, wire416, wire417, wire418, wire419, wire420, wire421, wire422, wire423, wire424, wire425, wire426, wire427, wire428, wire429, wire430, wire431, wire432, wire433, wire434, wire435, wire436, wire437, wire438, wire439, wire440, wire441, wire442, wire443, wire444, wire445, wire446, wire447, wire448, wire449, wire450, wire451, wire452, wire453, wire454, wire455, wire456, wire457, wire458, wire459, wire460, wire461, wire462, wire463, wire464, wire465, wire466, wire467, wire468, wire469, wire470, wire471, wire472, wire473, wire474, wire475, wire476, wire477, wire478, wire479, wire480, wire481, wire482, wire483, wire484, wire485, wire486, wire487, wire488, wire489, wire490, wire491, wire492, wire493, wire494, wire495, wire496, wire497, wire498, wire499, wire500, wire501, wire502, wire503, wire504, wire505, wire506, wire507, wire508, wire509, wire510, wire511, wire512, wire513, wire514, wire515, wire516, wire517, wire518, wire519, wire520, wire521, wire522, wire523, wire524, wire525, wire526, wire527, wire528, wire529, wire530, wire531, wire532, wire533, wire534, wire535, wire536, wire537, wire538, wire539, wire540, wire541, wire542, wire543, wire544, wire545, wire546, wire547, wire548, wire549, wire550, wire551, wire552, wire553, wire554, wire555, wire556, wire557, wire558, wire559, wire560, wire561, wire562, wire563, wire564, wire565, wire566, wire567, wire568, wire569, wire570, wire571, wire572, wire573, wire574, wire575, wire576, wire577, wire578, wire579, wire580, wire581, wire582, wire583, wire584, wire585, wire586, wire587, wire588, wire589, wire590, wire591, wire592, wire593, wire594, wire595, wire596, wire597, wire598, wire599, wire600, wire601, wire602, wire603, wire604, wire605, wire606, wire607, wire608, wire609, wire610, wire611, wire612, wire613, wire614, wire615, wire616, wire617, wire618, wire619, wire620, wire621, wire622, wire623, wire624, wire625, wire626, wire627, wire628, wire629, wire630, wire631, wire632, wire633, wire634, wire635, wire636, wire637, wire638, wire639, wire640, wire641, wire642, wire643, wire644, wire645, wire646, wire647, wire648, wire649, wire650, wire651, wire652, wire653, wire654, wire655, wire656, wire657, wire658, wire659, wire660, wire661, wire662, wire663, wire664, wire665, wire666, wire667, wire668, wire669, wire670, wire671, wire672, wire673, wire674, wire675, wire676, wire677, wire678, wire679, wire680, wire681, wire682, wire683, wire684, wire685, wire686, wire687, wire688, wire689, wire690, wire691, wire692, wire693, wire694, wire695, wire696, wire697, wire698, wire699, wire700, wire701, wire702, wire703, wire704, wire705, wire706, wire707, wire708, wire709, wire710, wire711, wire712, wire713, wire714, wire715, wire716, wire717, wire718, wire719, wire720, wire721, wire722, wire723, wire724, wire725, wire726, wire727, wire728, wire729, wire730, wire731, wire732, wire733, wire734, wire735, wire736, wire737, wire738, wire739, wire740, wire741, wire742, wire743, wire744, wire745, wire746, wire747, wire748, wire749, wire750, wire751, wire752, wire753, wire754, wire755, wire756, wire757, wire758, wire759, wire760, wire761, wire762, wire763, wire764, wire765, wire766, wire767, wire768, wire769, wire770, wire771, wire772, wire773, wire774, wire775, wire776, wire777, wire778, wire779, wire780, wire781, wire782, wire783, wire784, wire785, wire786, wire787, wire788, wire789, wire790, wire791, wire792, wire793, wire794, wire795, wire796, wire797, wire798, wire799, wire800, wire801, wire802, wire803, wire804, wire805, wire806, wire807, wire808, wire809, wire810, wire811, wire812, wire813, wire814, wire815, wire816, wire817, wire818, wire819, wire820, wire821, wire822, wire823, wire824, wire825, wire826, wire827, wire828, wire829, wire830, wire831, wire832, wire833, wire834, wire835, wire836, wire837, wire838, wire839, wire840, wire841, wire842, wire843, wire844, wire845, wire846, wire847, wire848, wire849, wire850, wire851, wire852, wire853, wire854, wire855, wire856, wire857, wire858, wire859, wire860, wire861, wire862, wire863, wire864, wire865, wire866, wire867, wire868, wire869, wire870, wire871, wire872, wire873, wire874, wire875, wire876, wire877, wire878, wire879, wire880, wire881, wire882, wire883, wire884, wire885, wire886, wire887, wire888, wire889, wire890, wire891, wire892, wire893, wire894, wire895, wire896, wire897, wire898, wire899, wire900, wire901, wire902, wire903, wire904, wire905, wire906, wire907, wire908, wire909, wire910, wire911, wire912, wire913, wire914, wire915, wire916, wire917, wire918, wire919, wire920, wire921, wire922, wire923, wire924, wire925, wire926, wire927, wire928, wire929, wire930, wire931, wire932, wire933, wire934, wire935, wire936, wire937, wire938, wire939, wire940, wire941, wire942, wire943, wire944, wire945, wire946, wire947, wire948, wire949, wire950, wire951, wire952, wire953, wire954, wire955, wire956, wire957, wire958, wire959, wire960, wire961, wire962, wire963, wire964, wire965, wire966, wire967, wire968, wire969, wire970, wire971, wire972, wire973, wire974, wire975, wire976, wire977, wire978, wire979, wire980, wire981, wire982, wire983, wire984, wire985, wire986, wire987, wire988, wire989, wire990, wire991, wire992, wire993, wire994, wire995, wire996, wire997, wire998, wire999, wire1000, wire1001, wire1002, wire1003, wire1004, wire1005, wire1006, wire1007, wire1008, wire1009, wire1010, wire1011, wire1012, wire1013, wire1014, wire1015, wire1016, wire1017, wire1018, wire1019, wire1020, wire1021, wire1022, wire1023, wire1024, wire1025, wire1026, wire1027, wire1028, wire1029, wire1030, wire1031, wire1032, wire1033, wire1034, wire1035, wire1036, wire1037, wire1038, wire1039, wire1040, wire1041, wire1042, wire1043, wire1044, wire1045, wire1046, wire1047, wire1048, wire1049, wire1050, wire1051, wire1052, wire1053, wire1054, wire1055, wire1056, wire1057, wire1058, wire1059, wire1060, wire1061, wire1062, wire1063, wire1064, wire1065, wire1066, wire1067, wire1068, wire1069, wire1070, wire1071, wire1072, wire1073, wire1074, wire1075, wire1076, wire1077, wire1078, wire1079, wire1080, wire1081, wire1082, wire1083, wire1084, wire1085, wire1086, wire1087, wire1088, wire1089, wire1090, wire1091, wire1092, wire1093, wire1094, wire1095, wire1096, wire1097, wire1098, wire1099, wire1100, wire1101, wire1102, wire1103, wire1104, wire1105, wire1106, wire1107, wire1108, wire1109, wire1110, wire1111, wire1112, wire1113, wire1114, wire1115, wire1116, wire1117, wire1118, wire1119, wire1120, wire1121, wire1122, wire1123, wire1124, wire1125, wire1126, wire1127, wire1128, wire1129, wire1130, wire1131, wire1132, wire1133, wire1134, wire1135, wire1136, wire1137, wire1138, wire1139, wire1140, wire1141, wire1142, wire1143, wire1144, wire1145, wire1146, wire1147, wire1148, wire1149, wire1150, wire1151, wire1152, wire1153, wire1154, wire1155, wire1156, wire1157, wire1158, wire1159, wire1160, wire1161, wire1162, wire1163, wire1164, wire1165, wire1166, wire1167, wire1168, wire1169, wire1170, wire1171, wire1172, wire1173, wire1174, wire1175, wire1176, wire1177, wire1178, wire1179, wire1180, wire1181, wire1182, wire1183, wire1184, wire1185, wire1186, wire1187, wire1188, wire1189, wire1190, wire1191, wire1192, wire1193, wire1194, wire1195, wire1196, wire1197, wire1198, wire1199, wire1200, wire1201, wire1202, wire1203, wire1204, wire1205, wire1206, wire1207, wire1208, wire1209, wire1210, wire1211, wire1212, wire1213, wire1214, wire1215, wire1216, wire1217, wire1218, wire1219, wire1220, wire1221, wire1222, wire1223, wire1224, wire1225, wire1226, wire1227, wire1228, wire1229, wire1230, wire1231, wire1232, wire1233, wire1234, wire1235, wire1236, wire1237, wire1238, wire1239, wire1240, wire1241, wire1242, wire1243, wire1244, wire1245, wire1246, wire1247, wire1248, wire1249, wire1250, wire1251, wire1252, wire1253, wire1254, wire1255, wire1256, wire1257, wire1258, wire1259, wire1260, wire1261, wire1262, wire1263, wire1264, wire1265, wire1266, wire1267, wire1268, wire1269, wire1270, wire1271, wire1272, wire1273, wire1274, wire1275, wire1276, wire1277, wire1278, wire1279, wire1280, wire1281, wire1282, wire1283, wire1284, wire1285, wire1286, wire1287, wire1288, wire1289, wire1290, wire1291, wire1292, wire1293, wire1294, wire1295, wire1296, wire1297, wire1298, wire1299, wire1300, wire1301, wire1302, wire1303, wire1304, wire1305, wire1306, wire1307, wire1308, wire1309, wire1310, wire1311, wire1312, wire1313, wire1314, wire1315, wire1316, wire1317, wire1318, wire1319, wire1320, wire1321, wire1322, wire1323, wire1324, wire1325, wire1326, wire1327, wire1328, wire1329, wire1330, wire1331, wire1332, wire1333, wire1334, wire1335, wire1336, wire1337, wire1338, wire1339, wire1340, wire1341, wire1342, wire1343, wire1344, wire1345, wire1346, wire1347, wire1348, wire1349, wire1350, wire1351, wire1352, wire1353, wire1354, wire1355, wire1356, wire1357, wire1358, wire1359, wire1360, wire1361, wire1362, wire1363, wire1364, wire1365, wire1366, wire1367, wire1368, wire1369, wire1370, wire1371, wire1372, wire1373, wire1374, wire1375, wire1376, wire1377, wire1378, wire1379, wire1380, wire1381, wire1382, wire1383, wire1384, wire1385, wire1386, wire1387, wire1388, wire1389, wire1390, wire1391, wire1392, wire1393, wire1394, wire1395, wire1396, wire1397, wire1398, wire1399, wire1400, wire1401, wire1402, wire1403, wire1404, wire1405, wire1406, wire1407, wire1408, wire1409, wire1410, wire1411, wire1412, wire1413, wire1414, wire1415, wire1416, wire1417, wire1418, wire1419, wire1420, wire1421, wire1422, wire1423, wire1424, wire1425, wire1426, wire1427, wire1428, wire1429, wire1430, wire1431, wire1432, wire1433, wire1434, wire1435, wire1436, wire1437, wire1438, wire1439, wire1440, wire1441, wire1442, wire1443, wire1444, wire1445, wire1446, wire1447, wire1448, wire1449, wire1450, wire1451, wire1452, wire1453, wire1454, wire1455, wire1456, wire1457, wire1458, wire1459, wire1460, wire1461, wire1462, wire1463, wire1464, wire1465, wire1466, wire1467, wire1468, wire1469, wire1470, wire1471, wire1472, wire1473, wire1474, wire1475, wire1476, wire1477, wire1478, wire1479, wire1480, wire1481, wire1482, wire1483, wire1484, wire1485, wire1486, wire1487, wire1488, wire1489, wire1490, wire1491, wire1492, wire1493, wire1494, wire1495, wire1496, wire1497, wire1498, wire1499, wire1500, wire1501, wire1502, wire1503, wire1504, wire1505, wire1506, wire1507, wire1508, wire1509, wire1510, wire1511, wire1512, wire1513, wire1514, wire1515, wire1516, wire1517, wire1518, wire1519, wire1520, wire1521, wire1522, wire1523, wire1524, wire1525, wire1526, wire1527, wire1528, wire1529, wire1530, wire1531, wire1532, wire1533, wire1534, wire1535, wire1536, wire1537, wire1538, wire1539, wire1540, wire1541, wire1542, wire1543, wire1544, wire1545, wire1546, wire1547, wire1548, wire1549, wire1550, wire1551, wire1552, wire1553, wire1554, wire1555, wire1556, wire1557, wire1558, wire1559, wire1560, wire1561, wire1562, wire1563, wire1564, wire1565, wire1566, wire1567, wire1568, wire1569, wire1570, wire1571, wire1572, wire1573, wire1574, wire1575, wire1576, wire1577, wire1578, wire1579, wire1580, wire1581, wire1582, wire1583, wire1584, wire1585, wire1586, wire1587, wire1588, wire1589, wire1590, wire1591, wire1592, wire1593, wire1594, wire1595, wire1596, wire1597, wire1598, wire1599, wire1600, wire1601, wire1602, wire1603, wire1604, wire1605, wire1606, wire1607, wire1608, wire1609, wire1610, wire1611, wire1612, wire1613, wire1614, wire1615, wire1616, wire1617, wire1618, wire1619, wire1620, wire1621, wire1622, wire1623, wire1624, wire1625, wire1626, wire1627, wire1628, wire1629, wire1630, wire1631, wire1632, wire1633, wire1634, wire1635, wire1636, wire1637, wire1638, wire1639, wire1640, wire1641, wire1642, wire1643, wire1644, wire1645, wire1646, wire1647, wire1648, wire1649, wire1650, wire1651, wire1652, wire1653, wire1654, wire1655, wire1656, wire1657, wire1658, wire1659, wire1660, wire1661, wire1662, wire1663, wire1664, wire1665, wire1666, wire1667, wire1668, wire1669, wire1670, wire1671, wire1672, wire1673, wire1674, wire1675, wire1676, wire1677, wire1678, wire1679, wire1680, wire1681, wire1682, wire1683, wire1684, wire1685, wire1686, wire1687, wire1688, wire1689, wire1690, wire1691, wire1692, wire1693, wire1694, wire1695, wire1696, wire1697, wire1698, wire1699, wire1700, wire1701, wire1702, wire1703, wire1704, wire1705, wire1706, wire1707, wire1708, wire1709, wire1710, wire1711, wire1712, wire1713, wire1714, wire1715, wire1716, wire1717, wire1718, wire1719, wire1720, wire1721, wire1722, wire1723, wire1724, wire1725, wire1726, wire1727, wire1728, wire1729, wire1730, wire1731, wire1732, wire1733, wire1734, wire1735, wire1736, wire1737, wire1738, wire1739, wire1740, wire1741, wire1742, wire1743, wire1744, wire1745, wire1746, wire1747, wire1748, wire1749, wire1750, wire1751, wire1752, wire1753, wire1754, wire1755, wire1756, wire1757, wire1758, wire1759, wire1760, wire1761, wire1762, wire1763, wire1764, wire1765, wire1766, wire1767, wire1768, wire1769, wire1770, wire1771, wire1772, wire1773, wire1774, wire1775, wire1776, wire1777, wire1778, wire1779, wire1780, wire1781, wire1782, wire1783, wire1784, wire1785, wire1786, wire1787, wire1788, wire1789, wire1790, wire1791, wire1792, wire1793, wire1794, wire1795, wire1796, wire1797, wire1798, wire1799, wire1800, wire1801, wire1802, wire1803, wire1804, wire1805, wire1806, wire1807, wire1808, wire1809, wire1810, wire1811, wire1812, wire1813, wire1814, wire1815, wire1816, wire1817, wire1818, wire1819, wire1820, wire1821, wire1822, wire1823, wire1824, wire1825, wire1826, wire1827, wire1828, wire1829, wire1830, wire1831, wire1832, wire1833, wire1834, wire1835, wire1836, wire1837, wire1838, wire1839, wire1840, wire1841, wire1842, wire1843, wire1844, wire1845, wire1846, wire1847, wire1848, wire1849, wire1850, wire1851, wire1852, wire1853, wire1854, wire1855, wire1856, wire1857, wire1858, wire1859, wire1860, wire1861, wire1862, wire1863, wire1864, wire1865, wire1866, wire1867, wire1868, wire1869, wire1870, wire1871, wire1872, wire1873, wire1874, wire1875, wire1876, wire1877, wire1878, wire1879, wire1880, wire1881, wire1882, wire1883, wire1884, wire1885, wire1886, wire1887, wire1888, wire1889, wire1890, wire1891, wire1892, wire1893, wire1894, wire1895, wire1896, wire1897, wire1898, wire1899, wire1900, wire1901, wire1902, wire1903, wire1904, wire1905, wire1906, wire1907, wire1908, wire1909, wire1910, wire1911, wire1912, wire1913, wire1914, wire1915, wire1916, wire1917, wire1918, wire1919, wire1920, wire1921, wire1922, wire1923, wire1924, wire1925, wire1926, wire1927, wire1928, wire1929, wire1930, wire1931, wire1932, wire1933, wire1934, wire1935, wire1936, wire1937, wire1938, wire1939, wire1940, wire1941, wire1942, wire1943, wire1944, wire1945, wire1946, wire1947, wire1948, wire1949, wire1950, wire1951, wire1952, wire1953, wire1954, wire1955, wire1956, wire1957, wire1958, wire1959, wire1960, wire1961, wire1962, wire1963, wire1964, wire1965, wire1966, wire1967, wire1968, wire1969, wire1970, wire1971, wire1972, wire1973, wire1974, wire1975, wire1976, wire1977, wire1978, wire1979, wire1980, wire1981, wire1982, wire1983, wire1984, wire1985, wire1986, wire1987, wire1988, wire1989, wire1990, wire1991, wire1992, wire1993, wire1994, wire1995, wire1996, wire1997, wire1998, wire1999, wire2000, wire2001, wire2002, wire2003, wire2004, wire2005, wire2006, wire2007, wire2008, wire2009, wire2010, wire2011, wire2012, wire2013, wire2014, wire2015, wire2016, wire2017, wire2018, wire2019, wire2020, wire2021, wire2022, wire2023, wire2024, wire2025, wire2026, wire2027, wire2028, wire2029, wire2030, wire2031, wire2032, wire2033, wire2034, wire2035, wire2036, wire2037, wire2038, wire2039, wire2040, wire2041, wire2042, wire2043, wire2044, wire2045, wire2046, wire2047, wire2048, wire2049, wire2050, wire2051, wire2052, wire2053, wire2054, wire2055, wire2056, wire2057, wire2058, wire2059, wire2060, wire2061, wire2062, wire2063, wire2064, wire2065, wire2066, wire2067, wire2068, wire2069, wire2070, wire2071, wire2072, wire2073, wire2074, wire2075, wire2076, wire2077, wire2078, wire2079, wire2080, wire2081, wire2082, wire2083, wire2084, wire2085, wire2086, wire2087, wire2088, wire2089, wire2090, wire2091, wire2092, wire2093, wire2094, wire2095, wire2096, wire2097, wire2098, wire2099, wire2100, wire2101, wire2102, wire2103, wire2104, wire2105, wire2106, wire2107, wire2108, wire2109, wire2110, wire2111, wire2112, wire2113, wire2114, wire2115, wire2116, wire2117, wire2118, wire2119, wire2120, wire2121, wire2122, wire2123, wire2124, wire2125, wire2126, wire2127, wire2128, wire2129, wire2130, wire2131, wire2132, wire2133, wire2134, wire2135, wire2136, wire2137, wire2138, wire2139, wire2140, wire2141, wire2142, wire2143, wire2144, wire2145, wire2146, wire2147, wire2148, wire2149, wire2150, wire2151, wire2152, wire2153, wire2154, wire2155, wire2156, wire2157, wire2158, wire2159, wire2160, wire2161, wire2162, wire2163, wire2164, wire2165, wire2166, wire2167, wire2168, wire2169, wire2170, wire2171, wire2172, wire2173, wire2174, wire2175, wire2176, wire2177, wire2178, wire2179, wire2180, wire2181, wire2182, wire2183, wire2184, wire2185, wire2186, wire2187, wire2188, wire2189, wire2190, wire2191, wire2192, wire2193, wire2194, wire2195, wire2196, wire2197, wire2198, wire2199, wire2200, wire2201, wire2202, wire2203, wire2204, wire2205, wire2206, wire2207, wire2208, wire2209, wire2210, wire2211, wire2212, wire2213, wire2214, wire2215, wire2216, wire2217, wire2218, wire2219, wire2220, wire2221, wire2222, wire2223, wire2224, wire2225, wire2226, wire2227, wire2228, wire2229, wire2230, wire2231, wire2232, wire2233, wire2234, wire2235, wire2236, wire2237, wire2238, wire2239, wire2240, wire2241, wire2242, wire2243, wire2244, wire2245, wire2246, wire2247, wire2248, wire2249, wire2250, wire2251, wire2252, wire2253, wire2254, wire2255, wire2256, wire2257, wire2258, wire2259, wire2260, wire2261, wire2262, wire2263, wire2264, wire2265, wire2266, wire2267, wire2268, wire2269, wire2270, wire2271, wire2272, wire2273, wire2274, wire2275, wire2276, wire2277, wire2278, wire2279, wire2280, wire2281, wire2282, wire2283, wire2284, wire2285, wire2286, wire2287, wire2288, wire2289, wire2290, wire2291, wire2292, wire2293, wire2294, wire2295, wire2296, wire2297, wire2298, wire2299, wire2300, wire2301, wire2302, wire2303, wire2304, wire2305, wire2306, wire2307, wire2308, wire2309, wire2310, wire2311, wire2312, wire2313, wire2314, wire2315, wire2316, wire2317, wire2318, wire2319, wire2320, wire2321, wire2322, wire2323, wire2324, wire2325, wire2326, wire2327, wire2328, wire2329, wire2330, wire2331, wire2332, wire2333, wire2334, wire2335, wire2336, wire2337, wire2338, wire2339, wire2340, wire2341, wire2342, wire2343, wire2344, wire2345, wire2346, wire2347, wire2348, wire2349, wire2350, wire2351, wire2352, wire2353, wire2354, wire2355, wire2356, wire2357, wire2358, wire2359, wire2360, wire2361, wire2362, wire2363, wire2364, wire2365, wire2366, wire2367, wire2368, wire2369, wire2370, wire2371, wire2372, wire2373, wire2374, wire2375, wire2376, wire2377, wire2378, wire2379, wire2380, wire2381, wire2382, wire2383, wire2384, wire2385, wire2386, wire2387, wire2388, wire2389, wire2390, wire2391, wire2392, wire2393, wire2394, wire2395, wire2396, wire2397, wire2398, wire2399, wire2400, wire2401, wire2402, wire2403, wire2404, wire2405, wire2406, wire2407, wire2408, wire2409, wire2410, wire2411, wire2412, wire2413, wire2414, wire2415, wire2416, wire2417, wire2418, wire2419, wire2420, wire2421, wire2422, wire2423, wire2424, wire2425, wire2426, wire2427, wire2428, wire2429, wire2430, wire2431, wire2432, wire2433, wire2434, wire2435, wire2436, wire2437, wire2438, wire2439, wire2440, wire2441, wire2442, wire2443, wire2444, wire2445, wire2446, wire2447, wire2448, wire2449, wire2450, wire2451, wire2452, wire2453, wire2454, wire2455, wire2456, wire2457, wire2458, wire2459, wire2460, wire2461, wire2462, wire2463, wire2464, wire2465, wire2466, wire2467, wire2468, wire2469, wire2470, wire2471, wire2472, wire2473, wire2474, wire2475, wire2476, wire2477, wire2478, wire2479, wire2480, wire2481, wire2482, wire2483, wire2484, wire2485, wire2486, wire2487, wire2488, wire2489, wire2490, wire2491, wire2492, wire2493, wire2494, wire2495, wire2496, wire2497, wire2498, wire2499, wire2500, wire2501, wire2502, wire2503, wire2504, wire2505, wire2506, wire2507, wire2508, wire2509, wire2510, wire2511, wire2512, wire2513, wire2514, wire2515, wire2516, wire2517, wire2518, wire2519, wire2520, wire2521, wire2522, wire2523, wire2524, wire2525, wire2526, wire2527, wire2528, wire2529, wire2530, wire2531, wire2532, wire2533, wire2534, wire2535, wire2536, wire2537, wire2538, wire2539, wire2540, wire2541, wire2542, wire2543, wire2544, wire2545, wire2546, wire2547, wire2548, wire2549, wire2550, wire2551, wire2552, wire2553, wire2554, wire2555, wire2556, wire2557, wire2558, wire2559, wire2560, wire2561, wire2562, wire2563, wire2564, wire2565, wire2566, wire2567, wire2568, wire2569, wire2570, wire2571, wire2572, wire2573, wire2574, wire2575, wire2576, wire2577, wire2578, wire2579, wire2580, wire2581, wire2582, wire2583, wire2584, wire2585, wire2586, wire2587, wire2588, wire2589, wire2590, wire2591, wire2592, wire2593, wire2594, wire2595, wire2596, wire2597, wire2598, wire2599, wire2600, wire2601, wire2602, wire2603, wire2604, wire2605, wire2606, wire2607, wire2608, wire2609, wire2610, wire2611, wire2612, wire2613, wire2614, wire2615, wire2616, wire2617, wire2618, wire2619, wire2620, wire2621, wire2622, wire2623, wire2624, wire2625, wire2626, wire2627, wire2628, wire2629, wire2630, wire2631, wire2632, wire2633, wire2634, wire2635, wire2636, wire2637, wire2638, wire2639, wire2640, wire2641, wire2642, wire2643, wire2644, wire2645, wire2646, wire2647, wire2648, wire2649, wire2650, wire2651, wire2652, wire2653, wire2654, wire2655, wire2656, wire2657, wire2658, wire2659, wire2660, wire2661, wire2662, wire2663, wire2664, wire2665, wire2666, wire2667, wire2668, wire2669, wire2670, wire2671, wire2672, wire2673, wire2674, wire2675, wire2676, wire2677, wire2678, wire2679, wire2680, wire2681, wire2682, wire2683, wire2684, wire2685, wire2686, wire2687, wire2688, wire2689, wire2690, wire2691, wire2692, wire2693, wire2694, wire2695, wire2696, wire2697, wire2698, wire2699, wire2700, wire2701, wire2702, wire2703, wire2704, wire2705, wire2706, wire2707, wire2708, wire2709, wire2710, wire2711, wire2712, wire2713, wire2714, wire2715, wire2716, wire2717, wire2718, wire2719, wire2720, wire2721, wire2722, wire2723, wire2724, wire2725, wire2726, wire2727, wire2728, wire2729, wire2730, wire2731, wire2732, wire2733, wire2734, wire2735, wire2736, wire2737, wire2738, wire2739, wire2740, wire2741, wire2742, wire2743, wire2744, wire2745, wire2746, wire2747, wire2748, wire2749, wire2750, wire2751, wire2752, wire2753, wire2754, wire2755, wire2756, wire2757, wire2758, wire2759, wire2760, wire2761, wire2762, wire2763, wire2764, wire2765, wire2766, wire2767, wire2768, wire2769, wire2770, wire2771, wire2772, wire2773, wire2774, wire2775, wire2776, wire2777, wire2778, wire2779, wire2780, wire2781, wire2782, wire2783, wire2784, wire2785, wire2786, wire2787, wire2788, wire2789, wire2790, wire2791, wire2792, wire2793, wire2794, wire2795, wire2796, wire2797, wire2798, wire2799, wire2800, wire2801, wire2802, wire2803, wire2804, wire2805, wire2806, wire2807, wire2808, wire2809, wire2810, wire2811, wire2812, wire2813, wire2814, wire2815, wire2816, wire2817, wire2818, wire2819, wire2820, wire2821, wire2822, wire2823, wire2824, wire2825, wire2826, wire2827, wire2828, wire2829, wire2830, wire2831, wire2832, wire2833, wire2834, wire2835, wire2836, wire2837, wire2838, wire2839, wire2840, wire2841, wire2842, wire2843, wire2844, wire2845, wire2846, wire2847, wire2848, wire2849, wire2850, wire2851, wire2852, wire2853, wire2854, wire2855, wire2856, wire2857, wire2858, wire2859, wire2860, wire2861, wire2862, wire2863, wire2864, wire2865, wire2866, wire2867, wire2868, wire2869, wire2870, wire2871, wire2872, wire2873, wire2874, wire2875, wire2876, wire2877, wire2878, wire2879, wire2880, wire2881, wire2882, wire2883, wire2884, wire2885, wire2886, wire2887, wire2888, wire2889, wire2890, wire2891, wire2892, wire2893, wire2894, wire2895, wire2896, wire2897, wire2898, wire2899, wire2900, wire2901, wire2902, wire2903, wire2904, wire2905, wire2906, wire2907, wire2908, wire2909, wire2910, wire2911, wire2912, wire2913, wire2914, wire2915, wire2916, wire2917, wire2918, wire2919, wire2920, wire2921, wire2922, wire2923, wire2924, wire2925, wire2926, wire2927, wire2928, wire2929, wire2930, wire2931, wire2932, wire2933, wire2934, wire2935, wire2936, wire2937, wire2938, wire2939, wire2940, wire2941, wire2942, wire2943, wire2944, wire2945, wire2946, wire2947, wire2948, wire2949, wire2950, wire2951, wire2952, wire2953, wire2954, wire2955, wire2956, wire2957, wire2958, wire2959, wire2960, wire2961, wire2962, wire2963, wire2964, wire2965, wire2966, wire2967, wire2968, wire2969, wire2970, wire2971, wire2972, wire2973, wire2974, wire2975, wire2976, wire2977, wire2978, wire2979, wire2980, wire2981, wire2982, wire2983, wire2984, wire2985, wire2986, wire2987, wire2988, wire2989, wire2990, wire2991, wire2992, wire2993, wire2994, wire2995, wire2996, wire2997, wire2998, wire2999, wire3000, wire3001, wire3002, wire3003, wire3004, wire3005, wire3006, wire3007, wire3008, wire3009, wire3010, wire3011, wire3012;

	and comp0(wire129, inA[0], inB[0]);
	and comp1(wire130, inA[0], inB[1]);
	and comp2(wire131, inA[0], inB[2]);
	and comp3(wire132, inA[0], inB[3]);
	and comp4(wire133, inA[0], inB[4]);
	and comp5(wire134, inA[0], inB[5]);
	and comp6(wire135, inA[0], inB[6]);
	and comp7(wire136, inA[0], inB[7]);
	and comp8(wire137, inA[0], inB[8]);
	and comp9(wire138, inA[0], inB[9]);
	and comp10(wire139, inA[0], inB[10]);
	and comp11(wire140, inA[0], inB[11]);
	and comp12(wire141, inA[0], inB[12]);
	and comp13(wire142, inA[0], inB[13]);
	and comp14(wire143, inA[0], inB[14]);
	and comp15(wire144, inA[0], inB[15]);
	and comp16(wire145, inA[0], inB[16]);
	and comp17(wire146, inA[0], inB[17]);
	and comp18(wire147, inA[0], inB[18]);
	and comp19(wire148, inA[0], inB[19]);
	and comp20(wire149, inA[0], inB[20]);
	and comp21(wire150, inA[0], inB[21]);
	and comp22(wire151, inA[0], inB[22]);
	and comp23(wire152, inA[0], inB[23]);
	and comp24(wire153, inA[0], inB[24]);
	and comp25(wire154, inA[0], inB[25]);
	and comp26(wire155, inA[0], inB[26]);
	and comp27(wire156, inA[0], inB[27]);
	and comp28(wire157, inA[0], inB[28]);
	and comp29(wire158, inA[0], inB[29]);
	and comp30(wire159, inA[0], inB[30]);
	and comp31(wire160, inA[0], inB[31]);
	and comp32(wire161, inA[1], inB[0]);
	and comp33(wire162, inA[1], inB[1]);
	and comp34(wire163, inA[1], inB[2]);
	and comp35(wire164, inA[1], inB[3]);
	and comp36(wire165, inA[1], inB[4]);
	and comp37(wire166, inA[1], inB[5]);
	and comp38(wire167, inA[1], inB[6]);
	and comp39(wire168, inA[1], inB[7]);
	and comp40(wire169, inA[1], inB[8]);
	and comp41(wire170, inA[1], inB[9]);
	and comp42(wire171, inA[1], inB[10]);
	and comp43(wire172, inA[1], inB[11]);
	and comp44(wire173, inA[1], inB[12]);
	and comp45(wire174, inA[1], inB[13]);
	and comp46(wire175, inA[1], inB[14]);
	and comp47(wire176, inA[1], inB[15]);
	and comp48(wire177, inA[1], inB[16]);
	and comp49(wire178, inA[1], inB[17]);
	and comp50(wire179, inA[1], inB[18]);
	and comp51(wire180, inA[1], inB[19]);
	and comp52(wire181, inA[1], inB[20]);
	and comp53(wire182, inA[1], inB[21]);
	and comp54(wire183, inA[1], inB[22]);
	and comp55(wire184, inA[1], inB[23]);
	and comp56(wire185, inA[1], inB[24]);
	and comp57(wire186, inA[1], inB[25]);
	and comp58(wire187, inA[1], inB[26]);
	and comp59(wire188, inA[1], inB[27]);
	and comp60(wire189, inA[1], inB[28]);
	and comp61(wire190, inA[1], inB[29]);
	and comp62(wire191, inA[1], inB[30]);
	and comp63(wire192, inA[1], inB[31]);
	and comp64(wire193, inA[2], inB[0]);
	and comp65(wire194, inA[2], inB[1]);
	and comp66(wire195, inA[2], inB[2]);
	and comp67(wire196, inA[2], inB[3]);
	and comp68(wire197, inA[2], inB[4]);
	and comp69(wire198, inA[2], inB[5]);
	and comp70(wire199, inA[2], inB[6]);
	and comp71(wire200, inA[2], inB[7]);
	and comp72(wire201, inA[2], inB[8]);
	and comp73(wire202, inA[2], inB[9]);
	and comp74(wire203, inA[2], inB[10]);
	and comp75(wire204, inA[2], inB[11]);
	and comp76(wire205, inA[2], inB[12]);
	and comp77(wire206, inA[2], inB[13]);
	and comp78(wire207, inA[2], inB[14]);
	and comp79(wire208, inA[2], inB[15]);
	and comp80(wire209, inA[2], inB[16]);
	and comp81(wire210, inA[2], inB[17]);
	and comp82(wire211, inA[2], inB[18]);
	and comp83(wire212, inA[2], inB[19]);
	and comp84(wire213, inA[2], inB[20]);
	and comp85(wire214, inA[2], inB[21]);
	and comp86(wire215, inA[2], inB[22]);
	and comp87(wire216, inA[2], inB[23]);
	and comp88(wire217, inA[2], inB[24]);
	and comp89(wire218, inA[2], inB[25]);
	and comp90(wire219, inA[2], inB[26]);
	and comp91(wire220, inA[2], inB[27]);
	and comp92(wire221, inA[2], inB[28]);
	and comp93(wire222, inA[2], inB[29]);
	and comp94(wire223, inA[2], inB[30]);
	and comp95(wire224, inA[2], inB[31]);
	and comp96(wire225, inA[3], inB[0]);
	and comp97(wire226, inA[3], inB[1]);
	and comp98(wire227, inA[3], inB[2]);
	and comp99(wire228, inA[3], inB[3]);
	and comp100(wire229, inA[3], inB[4]);
	and comp101(wire230, inA[3], inB[5]);
	and comp102(wire231, inA[3], inB[6]);
	and comp103(wire232, inA[3], inB[7]);
	and comp104(wire233, inA[3], inB[8]);
	and comp105(wire234, inA[3], inB[9]);
	and comp106(wire235, inA[3], inB[10]);
	and comp107(wire236, inA[3], inB[11]);
	and comp108(wire237, inA[3], inB[12]);
	and comp109(wire238, inA[3], inB[13]);
	and comp110(wire239, inA[3], inB[14]);
	and comp111(wire240, inA[3], inB[15]);
	and comp112(wire241, inA[3], inB[16]);
	and comp113(wire242, inA[3], inB[17]);
	and comp114(wire243, inA[3], inB[18]);
	and comp115(wire244, inA[3], inB[19]);
	and comp116(wire245, inA[3], inB[20]);
	and comp117(wire246, inA[3], inB[21]);
	and comp118(wire247, inA[3], inB[22]);
	and comp119(wire248, inA[3], inB[23]);
	and comp120(wire249, inA[3], inB[24]);
	and comp121(wire250, inA[3], inB[25]);
	and comp122(wire251, inA[3], inB[26]);
	and comp123(wire252, inA[3], inB[27]);
	and comp124(wire253, inA[3], inB[28]);
	and comp125(wire254, inA[3], inB[29]);
	and comp126(wire255, inA[3], inB[30]);
	and comp127(wire256, inA[3], inB[31]);
	and comp128(wire257, inA[4], inB[0]);
	and comp129(wire258, inA[4], inB[1]);
	and comp130(wire259, inA[4], inB[2]);
	and comp131(wire260, inA[4], inB[3]);
	and comp132(wire261, inA[4], inB[4]);
	and comp133(wire262, inA[4], inB[5]);
	and comp134(wire263, inA[4], inB[6]);
	and comp135(wire264, inA[4], inB[7]);
	and comp136(wire265, inA[4], inB[8]);
	and comp137(wire266, inA[4], inB[9]);
	and comp138(wire267, inA[4], inB[10]);
	and comp139(wire268, inA[4], inB[11]);
	and comp140(wire269, inA[4], inB[12]);
	and comp141(wire270, inA[4], inB[13]);
	and comp142(wire271, inA[4], inB[14]);
	and comp143(wire272, inA[4], inB[15]);
	and comp144(wire273, inA[4], inB[16]);
	and comp145(wire274, inA[4], inB[17]);
	and comp146(wire275, inA[4], inB[18]);
	and comp147(wire276, inA[4], inB[19]);
	and comp148(wire277, inA[4], inB[20]);
	and comp149(wire278, inA[4], inB[21]);
	and comp150(wire279, inA[4], inB[22]);
	and comp151(wire280, inA[4], inB[23]);
	and comp152(wire281, inA[4], inB[24]);
	and comp153(wire282, inA[4], inB[25]);
	and comp154(wire283, inA[4], inB[26]);
	and comp155(wire284, inA[4], inB[27]);
	and comp156(wire285, inA[4], inB[28]);
	and comp157(wire286, inA[4], inB[29]);
	and comp158(wire287, inA[4], inB[30]);
	and comp159(wire288, inA[4], inB[31]);
	and comp160(wire289, inA[5], inB[0]);
	and comp161(wire290, inA[5], inB[1]);
	and comp162(wire291, inA[5], inB[2]);
	and comp163(wire292, inA[5], inB[3]);
	and comp164(wire293, inA[5], inB[4]);
	and comp165(wire294, inA[5], inB[5]);
	and comp166(wire295, inA[5], inB[6]);
	and comp167(wire296, inA[5], inB[7]);
	and comp168(wire297, inA[5], inB[8]);
	and comp169(wire298, inA[5], inB[9]);
	and comp170(wire299, inA[5], inB[10]);
	and comp171(wire300, inA[5], inB[11]);
	and comp172(wire301, inA[5], inB[12]);
	and comp173(wire302, inA[5], inB[13]);
	and comp174(wire303, inA[5], inB[14]);
	and comp175(wire304, inA[5], inB[15]);
	and comp176(wire305, inA[5], inB[16]);
	and comp177(wire306, inA[5], inB[17]);
	and comp178(wire307, inA[5], inB[18]);
	and comp179(wire308, inA[5], inB[19]);
	and comp180(wire309, inA[5], inB[20]);
	and comp181(wire310, inA[5], inB[21]);
	and comp182(wire311, inA[5], inB[22]);
	and comp183(wire312, inA[5], inB[23]);
	and comp184(wire313, inA[5], inB[24]);
	and comp185(wire314, inA[5], inB[25]);
	and comp186(wire315, inA[5], inB[26]);
	and comp187(wire316, inA[5], inB[27]);
	and comp188(wire317, inA[5], inB[28]);
	and comp189(wire318, inA[5], inB[29]);
	and comp190(wire319, inA[5], inB[30]);
	and comp191(wire320, inA[5], inB[31]);
	and comp192(wire321, inA[6], inB[0]);
	and comp193(wire322, inA[6], inB[1]);
	and comp194(wire323, inA[6], inB[2]);
	and comp195(wire324, inA[6], inB[3]);
	and comp196(wire325, inA[6], inB[4]);
	and comp197(wire326, inA[6], inB[5]);
	and comp198(wire327, inA[6], inB[6]);
	and comp199(wire328, inA[6], inB[7]);
	and comp200(wire329, inA[6], inB[8]);
	and comp201(wire330, inA[6], inB[9]);
	and comp202(wire331, inA[6], inB[10]);
	and comp203(wire332, inA[6], inB[11]);
	and comp204(wire333, inA[6], inB[12]);
	and comp205(wire334, inA[6], inB[13]);
	and comp206(wire335, inA[6], inB[14]);
	and comp207(wire336, inA[6], inB[15]);
	and comp208(wire337, inA[6], inB[16]);
	and comp209(wire338, inA[6], inB[17]);
	and comp210(wire339, inA[6], inB[18]);
	and comp211(wire340, inA[6], inB[19]);
	and comp212(wire341, inA[6], inB[20]);
	and comp213(wire342, inA[6], inB[21]);
	and comp214(wire343, inA[6], inB[22]);
	and comp215(wire344, inA[6], inB[23]);
	and comp216(wire345, inA[6], inB[24]);
	and comp217(wire346, inA[6], inB[25]);
	and comp218(wire347, inA[6], inB[26]);
	and comp219(wire348, inA[6], inB[27]);
	and comp220(wire349, inA[6], inB[28]);
	and comp221(wire350, inA[6], inB[29]);
	and comp222(wire351, inA[6], inB[30]);
	and comp223(wire352, inA[6], inB[31]);
	and comp224(wire353, inA[7], inB[0]);
	and comp225(wire354, inA[7], inB[1]);
	and comp226(wire355, inA[7], inB[2]);
	and comp227(wire356, inA[7], inB[3]);
	and comp228(wire357, inA[7], inB[4]);
	and comp229(wire358, inA[7], inB[5]);
	and comp230(wire359, inA[7], inB[6]);
	and comp231(wire360, inA[7], inB[7]);
	and comp232(wire361, inA[7], inB[8]);
	and comp233(wire362, inA[7], inB[9]);
	and comp234(wire363, inA[7], inB[10]);
	and comp235(wire364, inA[7], inB[11]);
	and comp236(wire365, inA[7], inB[12]);
	and comp237(wire366, inA[7], inB[13]);
	and comp238(wire367, inA[7], inB[14]);
	and comp239(wire368, inA[7], inB[15]);
	and comp240(wire369, inA[7], inB[16]);
	and comp241(wire370, inA[7], inB[17]);
	and comp242(wire371, inA[7], inB[18]);
	and comp243(wire372, inA[7], inB[19]);
	and comp244(wire373, inA[7], inB[20]);
	and comp245(wire374, inA[7], inB[21]);
	and comp246(wire375, inA[7], inB[22]);
	and comp247(wire376, inA[7], inB[23]);
	and comp248(wire377, inA[7], inB[24]);
	and comp249(wire378, inA[7], inB[25]);
	and comp250(wire379, inA[7], inB[26]);
	and comp251(wire380, inA[7], inB[27]);
	and comp252(wire381, inA[7], inB[28]);
	and comp253(wire382, inA[7], inB[29]);
	and comp254(wire383, inA[7], inB[30]);
	and comp255(wire384, inA[7], inB[31]);
	and comp256(wire385, inA[8], inB[0]);
	and comp257(wire386, inA[8], inB[1]);
	and comp258(wire387, inA[8], inB[2]);
	and comp259(wire388, inA[8], inB[3]);
	and comp260(wire389, inA[8], inB[4]);
	and comp261(wire390, inA[8], inB[5]);
	and comp262(wire391, inA[8], inB[6]);
	and comp263(wire392, inA[8], inB[7]);
	and comp264(wire393, inA[8], inB[8]);
	and comp265(wire394, inA[8], inB[9]);
	and comp266(wire395, inA[8], inB[10]);
	and comp267(wire396, inA[8], inB[11]);
	and comp268(wire397, inA[8], inB[12]);
	and comp269(wire398, inA[8], inB[13]);
	and comp270(wire399, inA[8], inB[14]);
	and comp271(wire400, inA[8], inB[15]);
	and comp272(wire401, inA[8], inB[16]);
	and comp273(wire402, inA[8], inB[17]);
	and comp274(wire403, inA[8], inB[18]);
	and comp275(wire404, inA[8], inB[19]);
	and comp276(wire405, inA[8], inB[20]);
	and comp277(wire406, inA[8], inB[21]);
	and comp278(wire407, inA[8], inB[22]);
	and comp279(wire408, inA[8], inB[23]);
	and comp280(wire409, inA[8], inB[24]);
	and comp281(wire410, inA[8], inB[25]);
	and comp282(wire411, inA[8], inB[26]);
	and comp283(wire412, inA[8], inB[27]);
	and comp284(wire413, inA[8], inB[28]);
	and comp285(wire414, inA[8], inB[29]);
	and comp286(wire415, inA[8], inB[30]);
	and comp287(wire416, inA[8], inB[31]);
	and comp288(wire417, inA[9], inB[0]);
	and comp289(wire418, inA[9], inB[1]);
	and comp290(wire419, inA[9], inB[2]);
	and comp291(wire420, inA[9], inB[3]);
	and comp292(wire421, inA[9], inB[4]);
	and comp293(wire422, inA[9], inB[5]);
	and comp294(wire423, inA[9], inB[6]);
	and comp295(wire424, inA[9], inB[7]);
	and comp296(wire425, inA[9], inB[8]);
	and comp297(wire426, inA[9], inB[9]);
	and comp298(wire427, inA[9], inB[10]);
	and comp299(wire428, inA[9], inB[11]);
	and comp300(wire429, inA[9], inB[12]);
	and comp301(wire430, inA[9], inB[13]);
	and comp302(wire431, inA[9], inB[14]);
	and comp303(wire432, inA[9], inB[15]);
	and comp304(wire433, inA[9], inB[16]);
	and comp305(wire434, inA[9], inB[17]);
	and comp306(wire435, inA[9], inB[18]);
	and comp307(wire436, inA[9], inB[19]);
	and comp308(wire437, inA[9], inB[20]);
	and comp309(wire438, inA[9], inB[21]);
	and comp310(wire439, inA[9], inB[22]);
	and comp311(wire440, inA[9], inB[23]);
	and comp312(wire441, inA[9], inB[24]);
	and comp313(wire442, inA[9], inB[25]);
	and comp314(wire443, inA[9], inB[26]);
	and comp315(wire444, inA[9], inB[27]);
	and comp316(wire445, inA[9], inB[28]);
	and comp317(wire446, inA[9], inB[29]);
	and comp318(wire447, inA[9], inB[30]);
	and comp319(wire448, inA[9], inB[31]);
	and comp320(wire449, inA[10], inB[0]);
	and comp321(wire450, inA[10], inB[1]);
	and comp322(wire451, inA[10], inB[2]);
	and comp323(wire452, inA[10], inB[3]);
	and comp324(wire453, inA[10], inB[4]);
	and comp325(wire454, inA[10], inB[5]);
	and comp326(wire455, inA[10], inB[6]);
	and comp327(wire456, inA[10], inB[7]);
	and comp328(wire457, inA[10], inB[8]);
	and comp329(wire458, inA[10], inB[9]);
	and comp330(wire459, inA[10], inB[10]);
	and comp331(wire460, inA[10], inB[11]);
	and comp332(wire461, inA[10], inB[12]);
	and comp333(wire462, inA[10], inB[13]);
	and comp334(wire463, inA[10], inB[14]);
	and comp335(wire464, inA[10], inB[15]);
	and comp336(wire465, inA[10], inB[16]);
	and comp337(wire466, inA[10], inB[17]);
	and comp338(wire467, inA[10], inB[18]);
	and comp339(wire468, inA[10], inB[19]);
	and comp340(wire469, inA[10], inB[20]);
	and comp341(wire470, inA[10], inB[21]);
	and comp342(wire471, inA[10], inB[22]);
	and comp343(wire472, inA[10], inB[23]);
	and comp344(wire473, inA[10], inB[24]);
	and comp345(wire474, inA[10], inB[25]);
	and comp346(wire475, inA[10], inB[26]);
	and comp347(wire476, inA[10], inB[27]);
	and comp348(wire477, inA[10], inB[28]);
	and comp349(wire478, inA[10], inB[29]);
	and comp350(wire479, inA[10], inB[30]);
	and comp351(wire480, inA[10], inB[31]);
	and comp352(wire481, inA[11], inB[0]);
	and comp353(wire482, inA[11], inB[1]);
	and comp354(wire483, inA[11], inB[2]);
	and comp355(wire484, inA[11], inB[3]);
	and comp356(wire485, inA[11], inB[4]);
	and comp357(wire486, inA[11], inB[5]);
	and comp358(wire487, inA[11], inB[6]);
	and comp359(wire488, inA[11], inB[7]);
	and comp360(wire489, inA[11], inB[8]);
	and comp361(wire490, inA[11], inB[9]);
	and comp362(wire491, inA[11], inB[10]);
	and comp363(wire492, inA[11], inB[11]);
	and comp364(wire493, inA[11], inB[12]);
	and comp365(wire494, inA[11], inB[13]);
	and comp366(wire495, inA[11], inB[14]);
	and comp367(wire496, inA[11], inB[15]);
	and comp368(wire497, inA[11], inB[16]);
	and comp369(wire498, inA[11], inB[17]);
	and comp370(wire499, inA[11], inB[18]);
	and comp371(wire500, inA[11], inB[19]);
	and comp372(wire501, inA[11], inB[20]);
	and comp373(wire502, inA[11], inB[21]);
	and comp374(wire503, inA[11], inB[22]);
	and comp375(wire504, inA[11], inB[23]);
	and comp376(wire505, inA[11], inB[24]);
	and comp377(wire506, inA[11], inB[25]);
	and comp378(wire507, inA[11], inB[26]);
	and comp379(wire508, inA[11], inB[27]);
	and comp380(wire509, inA[11], inB[28]);
	and comp381(wire510, inA[11], inB[29]);
	and comp382(wire511, inA[11], inB[30]);
	and comp383(wire512, inA[11], inB[31]);
	and comp384(wire513, inA[12], inB[0]);
	and comp385(wire514, inA[12], inB[1]);
	and comp386(wire515, inA[12], inB[2]);
	and comp387(wire516, inA[12], inB[3]);
	and comp388(wire517, inA[12], inB[4]);
	and comp389(wire518, inA[12], inB[5]);
	and comp390(wire519, inA[12], inB[6]);
	and comp391(wire520, inA[12], inB[7]);
	and comp392(wire521, inA[12], inB[8]);
	and comp393(wire522, inA[12], inB[9]);
	and comp394(wire523, inA[12], inB[10]);
	and comp395(wire524, inA[12], inB[11]);
	and comp396(wire525, inA[12], inB[12]);
	and comp397(wire526, inA[12], inB[13]);
	and comp398(wire527, inA[12], inB[14]);
	and comp399(wire528, inA[12], inB[15]);
	and comp400(wire529, inA[12], inB[16]);
	and comp401(wire530, inA[12], inB[17]);
	and comp402(wire531, inA[12], inB[18]);
	and comp403(wire532, inA[12], inB[19]);
	and comp404(wire533, inA[12], inB[20]);
	and comp405(wire534, inA[12], inB[21]);
	and comp406(wire535, inA[12], inB[22]);
	and comp407(wire536, inA[12], inB[23]);
	and comp408(wire537, inA[12], inB[24]);
	and comp409(wire538, inA[12], inB[25]);
	and comp410(wire539, inA[12], inB[26]);
	and comp411(wire540, inA[12], inB[27]);
	and comp412(wire541, inA[12], inB[28]);
	and comp413(wire542, inA[12], inB[29]);
	and comp414(wire543, inA[12], inB[30]);
	and comp415(wire544, inA[12], inB[31]);
	and comp416(wire545, inA[13], inB[0]);
	and comp417(wire546, inA[13], inB[1]);
	and comp418(wire547, inA[13], inB[2]);
	and comp419(wire548, inA[13], inB[3]);
	and comp420(wire549, inA[13], inB[4]);
	and comp421(wire550, inA[13], inB[5]);
	and comp422(wire551, inA[13], inB[6]);
	and comp423(wire552, inA[13], inB[7]);
	and comp424(wire553, inA[13], inB[8]);
	and comp425(wire554, inA[13], inB[9]);
	and comp426(wire555, inA[13], inB[10]);
	and comp427(wire556, inA[13], inB[11]);
	and comp428(wire557, inA[13], inB[12]);
	and comp429(wire558, inA[13], inB[13]);
	and comp430(wire559, inA[13], inB[14]);
	and comp431(wire560, inA[13], inB[15]);
	and comp432(wire561, inA[13], inB[16]);
	and comp433(wire562, inA[13], inB[17]);
	and comp434(wire563, inA[13], inB[18]);
	and comp435(wire564, inA[13], inB[19]);
	and comp436(wire565, inA[13], inB[20]);
	and comp437(wire566, inA[13], inB[21]);
	and comp438(wire567, inA[13], inB[22]);
	and comp439(wire568, inA[13], inB[23]);
	and comp440(wire569, inA[13], inB[24]);
	and comp441(wire570, inA[13], inB[25]);
	and comp442(wire571, inA[13], inB[26]);
	and comp443(wire572, inA[13], inB[27]);
	and comp444(wire573, inA[13], inB[28]);
	and comp445(wire574, inA[13], inB[29]);
	and comp446(wire575, inA[13], inB[30]);
	and comp447(wire576, inA[13], inB[31]);
	and comp448(wire577, inA[14], inB[0]);
	and comp449(wire578, inA[14], inB[1]);
	and comp450(wire579, inA[14], inB[2]);
	and comp451(wire580, inA[14], inB[3]);
	and comp452(wire581, inA[14], inB[4]);
	and comp453(wire582, inA[14], inB[5]);
	and comp454(wire583, inA[14], inB[6]);
	and comp455(wire584, inA[14], inB[7]);
	and comp456(wire585, inA[14], inB[8]);
	and comp457(wire586, inA[14], inB[9]);
	and comp458(wire587, inA[14], inB[10]);
	and comp459(wire588, inA[14], inB[11]);
	and comp460(wire589, inA[14], inB[12]);
	and comp461(wire590, inA[14], inB[13]);
	and comp462(wire591, inA[14], inB[14]);
	and comp463(wire592, inA[14], inB[15]);
	and comp464(wire593, inA[14], inB[16]);
	and comp465(wire594, inA[14], inB[17]);
	and comp466(wire595, inA[14], inB[18]);
	and comp467(wire596, inA[14], inB[19]);
	and comp468(wire597, inA[14], inB[20]);
	and comp469(wire598, inA[14], inB[21]);
	and comp470(wire599, inA[14], inB[22]);
	and comp471(wire600, inA[14], inB[23]);
	and comp472(wire601, inA[14], inB[24]);
	and comp473(wire602, inA[14], inB[25]);
	and comp474(wire603, inA[14], inB[26]);
	and comp475(wire604, inA[14], inB[27]);
	and comp476(wire605, inA[14], inB[28]);
	and comp477(wire606, inA[14], inB[29]);
	and comp478(wire607, inA[14], inB[30]);
	and comp479(wire608, inA[14], inB[31]);
	and comp480(wire609, inA[15], inB[0]);
	and comp481(wire610, inA[15], inB[1]);
	and comp482(wire611, inA[15], inB[2]);
	and comp483(wire612, inA[15], inB[3]);
	and comp484(wire613, inA[15], inB[4]);
	and comp485(wire614, inA[15], inB[5]);
	and comp486(wire615, inA[15], inB[6]);
	and comp487(wire616, inA[15], inB[7]);
	and comp488(wire617, inA[15], inB[8]);
	and comp489(wire618, inA[15], inB[9]);
	and comp490(wire619, inA[15], inB[10]);
	and comp491(wire620, inA[15], inB[11]);
	and comp492(wire621, inA[15], inB[12]);
	and comp493(wire622, inA[15], inB[13]);
	and comp494(wire623, inA[15], inB[14]);
	and comp495(wire624, inA[15], inB[15]);
	and comp496(wire625, inA[15], inB[16]);
	and comp497(wire626, inA[15], inB[17]);
	and comp498(wire627, inA[15], inB[18]);
	and comp499(wire628, inA[15], inB[19]);
	and comp500(wire629, inA[15], inB[20]);
	and comp501(wire630, inA[15], inB[21]);
	and comp502(wire631, inA[15], inB[22]);
	and comp503(wire632, inA[15], inB[23]);
	and comp504(wire633, inA[15], inB[24]);
	and comp505(wire634, inA[15], inB[25]);
	and comp506(wire635, inA[15], inB[26]);
	and comp507(wire636, inA[15], inB[27]);
	and comp508(wire637, inA[15], inB[28]);
	and comp509(wire638, inA[15], inB[29]);
	and comp510(wire639, inA[15], inB[30]);
	and comp511(wire640, inA[15], inB[31]);
	and comp512(wire641, inA[16], inB[0]);
	and comp513(wire642, inA[16], inB[1]);
	and comp514(wire643, inA[16], inB[2]);
	and comp515(wire644, inA[16], inB[3]);
	and comp516(wire645, inA[16], inB[4]);
	and comp517(wire646, inA[16], inB[5]);
	and comp518(wire647, inA[16], inB[6]);
	and comp519(wire648, inA[16], inB[7]);
	and comp520(wire649, inA[16], inB[8]);
	and comp521(wire650, inA[16], inB[9]);
	and comp522(wire651, inA[16], inB[10]);
	and comp523(wire652, inA[16], inB[11]);
	and comp524(wire653, inA[16], inB[12]);
	and comp525(wire654, inA[16], inB[13]);
	and comp526(wire655, inA[16], inB[14]);
	and comp527(wire656, inA[16], inB[15]);
	and comp528(wire657, inA[16], inB[16]);
	and comp529(wire658, inA[16], inB[17]);
	and comp530(wire659, inA[16], inB[18]);
	and comp531(wire660, inA[16], inB[19]);
	and comp532(wire661, inA[16], inB[20]);
	and comp533(wire662, inA[16], inB[21]);
	and comp534(wire663, inA[16], inB[22]);
	and comp535(wire664, inA[16], inB[23]);
	and comp536(wire665, inA[16], inB[24]);
	and comp537(wire666, inA[16], inB[25]);
	and comp538(wire667, inA[16], inB[26]);
	and comp539(wire668, inA[16], inB[27]);
	and comp540(wire669, inA[16], inB[28]);
	and comp541(wire670, inA[16], inB[29]);
	and comp542(wire671, inA[16], inB[30]);
	and comp543(wire672, inA[16], inB[31]);
	and comp544(wire673, inA[17], inB[0]);
	and comp545(wire674, inA[17], inB[1]);
	and comp546(wire675, inA[17], inB[2]);
	and comp547(wire676, inA[17], inB[3]);
	and comp548(wire677, inA[17], inB[4]);
	and comp549(wire678, inA[17], inB[5]);
	and comp550(wire679, inA[17], inB[6]);
	and comp551(wire680, inA[17], inB[7]);
	and comp552(wire681, inA[17], inB[8]);
	and comp553(wire682, inA[17], inB[9]);
	and comp554(wire683, inA[17], inB[10]);
	and comp555(wire684, inA[17], inB[11]);
	and comp556(wire685, inA[17], inB[12]);
	and comp557(wire686, inA[17], inB[13]);
	and comp558(wire687, inA[17], inB[14]);
	and comp559(wire688, inA[17], inB[15]);
	and comp560(wire689, inA[17], inB[16]);
	and comp561(wire690, inA[17], inB[17]);
	and comp562(wire691, inA[17], inB[18]);
	and comp563(wire692, inA[17], inB[19]);
	and comp564(wire693, inA[17], inB[20]);
	and comp565(wire694, inA[17], inB[21]);
	and comp566(wire695, inA[17], inB[22]);
	and comp567(wire696, inA[17], inB[23]);
	and comp568(wire697, inA[17], inB[24]);
	and comp569(wire698, inA[17], inB[25]);
	and comp570(wire699, inA[17], inB[26]);
	and comp571(wire700, inA[17], inB[27]);
	and comp572(wire701, inA[17], inB[28]);
	and comp573(wire702, inA[17], inB[29]);
	and comp574(wire703, inA[17], inB[30]);
	and comp575(wire704, inA[17], inB[31]);
	and comp576(wire705, inA[18], inB[0]);
	and comp577(wire706, inA[18], inB[1]);
	and comp578(wire707, inA[18], inB[2]);
	and comp579(wire708, inA[18], inB[3]);
	and comp580(wire709, inA[18], inB[4]);
	and comp581(wire710, inA[18], inB[5]);
	and comp582(wire711, inA[18], inB[6]);
	and comp583(wire712, inA[18], inB[7]);
	and comp584(wire713, inA[18], inB[8]);
	and comp585(wire714, inA[18], inB[9]);
	and comp586(wire715, inA[18], inB[10]);
	and comp587(wire716, inA[18], inB[11]);
	and comp588(wire717, inA[18], inB[12]);
	and comp589(wire718, inA[18], inB[13]);
	and comp590(wire719, inA[18], inB[14]);
	and comp591(wire720, inA[18], inB[15]);
	and comp592(wire721, inA[18], inB[16]);
	and comp593(wire722, inA[18], inB[17]);
	and comp594(wire723, inA[18], inB[18]);
	and comp595(wire724, inA[18], inB[19]);
	and comp596(wire725, inA[18], inB[20]);
	and comp597(wire726, inA[18], inB[21]);
	and comp598(wire727, inA[18], inB[22]);
	and comp599(wire728, inA[18], inB[23]);
	and comp600(wire729, inA[18], inB[24]);
	and comp601(wire730, inA[18], inB[25]);
	and comp602(wire731, inA[18], inB[26]);
	and comp603(wire732, inA[18], inB[27]);
	and comp604(wire733, inA[18], inB[28]);
	and comp605(wire734, inA[18], inB[29]);
	and comp606(wire735, inA[18], inB[30]);
	and comp607(wire736, inA[18], inB[31]);
	and comp608(wire737, inA[19], inB[0]);
	and comp609(wire738, inA[19], inB[1]);
	and comp610(wire739, inA[19], inB[2]);
	and comp611(wire740, inA[19], inB[3]);
	and comp612(wire741, inA[19], inB[4]);
	and comp613(wire742, inA[19], inB[5]);
	and comp614(wire743, inA[19], inB[6]);
	and comp615(wire744, inA[19], inB[7]);
	and comp616(wire745, inA[19], inB[8]);
	and comp617(wire746, inA[19], inB[9]);
	and comp618(wire747, inA[19], inB[10]);
	and comp619(wire748, inA[19], inB[11]);
	and comp620(wire749, inA[19], inB[12]);
	and comp621(wire750, inA[19], inB[13]);
	and comp622(wire751, inA[19], inB[14]);
	and comp623(wire752, inA[19], inB[15]);
	and comp624(wire753, inA[19], inB[16]);
	and comp625(wire754, inA[19], inB[17]);
	and comp626(wire755, inA[19], inB[18]);
	and comp627(wire756, inA[19], inB[19]);
	and comp628(wire757, inA[19], inB[20]);
	and comp629(wire758, inA[19], inB[21]);
	and comp630(wire759, inA[19], inB[22]);
	and comp631(wire760, inA[19], inB[23]);
	and comp632(wire761, inA[19], inB[24]);
	and comp633(wire762, inA[19], inB[25]);
	and comp634(wire763, inA[19], inB[26]);
	and comp635(wire764, inA[19], inB[27]);
	and comp636(wire765, inA[19], inB[28]);
	and comp637(wire766, inA[19], inB[29]);
	and comp638(wire767, inA[19], inB[30]);
	and comp639(wire768, inA[19], inB[31]);
	and comp640(wire769, inA[20], inB[0]);
	and comp641(wire770, inA[20], inB[1]);
	and comp642(wire771, inA[20], inB[2]);
	and comp643(wire772, inA[20], inB[3]);
	and comp644(wire773, inA[20], inB[4]);
	and comp645(wire774, inA[20], inB[5]);
	and comp646(wire775, inA[20], inB[6]);
	and comp647(wire776, inA[20], inB[7]);
	and comp648(wire777, inA[20], inB[8]);
	and comp649(wire778, inA[20], inB[9]);
	and comp650(wire779, inA[20], inB[10]);
	and comp651(wire780, inA[20], inB[11]);
	and comp652(wire781, inA[20], inB[12]);
	and comp653(wire782, inA[20], inB[13]);
	and comp654(wire783, inA[20], inB[14]);
	and comp655(wire784, inA[20], inB[15]);
	and comp656(wire785, inA[20], inB[16]);
	and comp657(wire786, inA[20], inB[17]);
	and comp658(wire787, inA[20], inB[18]);
	and comp659(wire788, inA[20], inB[19]);
	and comp660(wire789, inA[20], inB[20]);
	and comp661(wire790, inA[20], inB[21]);
	and comp662(wire791, inA[20], inB[22]);
	and comp663(wire792, inA[20], inB[23]);
	and comp664(wire793, inA[20], inB[24]);
	and comp665(wire794, inA[20], inB[25]);
	and comp666(wire795, inA[20], inB[26]);
	and comp667(wire796, inA[20], inB[27]);
	and comp668(wire797, inA[20], inB[28]);
	and comp669(wire798, inA[20], inB[29]);
	and comp670(wire799, inA[20], inB[30]);
	and comp671(wire800, inA[20], inB[31]);
	and comp672(wire801, inA[21], inB[0]);
	and comp673(wire802, inA[21], inB[1]);
	and comp674(wire803, inA[21], inB[2]);
	and comp675(wire804, inA[21], inB[3]);
	and comp676(wire805, inA[21], inB[4]);
	and comp677(wire806, inA[21], inB[5]);
	and comp678(wire807, inA[21], inB[6]);
	and comp679(wire808, inA[21], inB[7]);
	and comp680(wire809, inA[21], inB[8]);
	and comp681(wire810, inA[21], inB[9]);
	and comp682(wire811, inA[21], inB[10]);
	and comp683(wire812, inA[21], inB[11]);
	and comp684(wire813, inA[21], inB[12]);
	and comp685(wire814, inA[21], inB[13]);
	and comp686(wire815, inA[21], inB[14]);
	and comp687(wire816, inA[21], inB[15]);
	and comp688(wire817, inA[21], inB[16]);
	and comp689(wire818, inA[21], inB[17]);
	and comp690(wire819, inA[21], inB[18]);
	and comp691(wire820, inA[21], inB[19]);
	and comp692(wire821, inA[21], inB[20]);
	and comp693(wire822, inA[21], inB[21]);
	and comp694(wire823, inA[21], inB[22]);
	and comp695(wire824, inA[21], inB[23]);
	and comp696(wire825, inA[21], inB[24]);
	and comp697(wire826, inA[21], inB[25]);
	and comp698(wire827, inA[21], inB[26]);
	and comp699(wire828, inA[21], inB[27]);
	and comp700(wire829, inA[21], inB[28]);
	and comp701(wire830, inA[21], inB[29]);
	and comp702(wire831, inA[21], inB[30]);
	and comp703(wire832, inA[21], inB[31]);
	and comp704(wire833, inA[22], inB[0]);
	and comp705(wire834, inA[22], inB[1]);
	and comp706(wire835, inA[22], inB[2]);
	and comp707(wire836, inA[22], inB[3]);
	and comp708(wire837, inA[22], inB[4]);
	and comp709(wire838, inA[22], inB[5]);
	and comp710(wire839, inA[22], inB[6]);
	and comp711(wire840, inA[22], inB[7]);
	and comp712(wire841, inA[22], inB[8]);
	and comp713(wire842, inA[22], inB[9]);
	and comp714(wire843, inA[22], inB[10]);
	and comp715(wire844, inA[22], inB[11]);
	and comp716(wire845, inA[22], inB[12]);
	and comp717(wire846, inA[22], inB[13]);
	and comp718(wire847, inA[22], inB[14]);
	and comp719(wire848, inA[22], inB[15]);
	and comp720(wire849, inA[22], inB[16]);
	and comp721(wire850, inA[22], inB[17]);
	and comp722(wire851, inA[22], inB[18]);
	and comp723(wire852, inA[22], inB[19]);
	and comp724(wire853, inA[22], inB[20]);
	and comp725(wire854, inA[22], inB[21]);
	and comp726(wire855, inA[22], inB[22]);
	and comp727(wire856, inA[22], inB[23]);
	and comp728(wire857, inA[22], inB[24]);
	and comp729(wire858, inA[22], inB[25]);
	and comp730(wire859, inA[22], inB[26]);
	and comp731(wire860, inA[22], inB[27]);
	and comp732(wire861, inA[22], inB[28]);
	and comp733(wire862, inA[22], inB[29]);
	and comp734(wire863, inA[22], inB[30]);
	and comp735(wire864, inA[22], inB[31]);
	and comp736(wire865, inA[23], inB[0]);
	and comp737(wire866, inA[23], inB[1]);
	and comp738(wire867, inA[23], inB[2]);
	and comp739(wire868, inA[23], inB[3]);
	and comp740(wire869, inA[23], inB[4]);
	and comp741(wire870, inA[23], inB[5]);
	and comp742(wire871, inA[23], inB[6]);
	and comp743(wire872, inA[23], inB[7]);
	and comp744(wire873, inA[23], inB[8]);
	and comp745(wire874, inA[23], inB[9]);
	and comp746(wire875, inA[23], inB[10]);
	and comp747(wire876, inA[23], inB[11]);
	and comp748(wire877, inA[23], inB[12]);
	and comp749(wire878, inA[23], inB[13]);
	and comp750(wire879, inA[23], inB[14]);
	and comp751(wire880, inA[23], inB[15]);
	and comp752(wire881, inA[23], inB[16]);
	and comp753(wire882, inA[23], inB[17]);
	and comp754(wire883, inA[23], inB[18]);
	and comp755(wire884, inA[23], inB[19]);
	and comp756(wire885, inA[23], inB[20]);
	and comp757(wire886, inA[23], inB[21]);
	and comp758(wire887, inA[23], inB[22]);
	and comp759(wire888, inA[23], inB[23]);
	and comp760(wire889, inA[23], inB[24]);
	and comp761(wire890, inA[23], inB[25]);
	and comp762(wire891, inA[23], inB[26]);
	and comp763(wire892, inA[23], inB[27]);
	and comp764(wire893, inA[23], inB[28]);
	and comp765(wire894, inA[23], inB[29]);
	and comp766(wire895, inA[23], inB[30]);
	and comp767(wire896, inA[23], inB[31]);
	and comp768(wire897, inA[24], inB[0]);
	and comp769(wire898, inA[24], inB[1]);
	and comp770(wire899, inA[24], inB[2]);
	and comp771(wire900, inA[24], inB[3]);
	and comp772(wire901, inA[24], inB[4]);
	and comp773(wire902, inA[24], inB[5]);
	and comp774(wire903, inA[24], inB[6]);
	and comp775(wire904, inA[24], inB[7]);
	and comp776(wire905, inA[24], inB[8]);
	and comp777(wire906, inA[24], inB[9]);
	and comp778(wire907, inA[24], inB[10]);
	and comp779(wire908, inA[24], inB[11]);
	and comp780(wire909, inA[24], inB[12]);
	and comp781(wire910, inA[24], inB[13]);
	and comp782(wire911, inA[24], inB[14]);
	and comp783(wire912, inA[24], inB[15]);
	and comp784(wire913, inA[24], inB[16]);
	and comp785(wire914, inA[24], inB[17]);
	and comp786(wire915, inA[24], inB[18]);
	and comp787(wire916, inA[24], inB[19]);
	and comp788(wire917, inA[24], inB[20]);
	and comp789(wire918, inA[24], inB[21]);
	and comp790(wire919, inA[24], inB[22]);
	and comp791(wire920, inA[24], inB[23]);
	and comp792(wire921, inA[24], inB[24]);
	and comp793(wire922, inA[24], inB[25]);
	and comp794(wire923, inA[24], inB[26]);
	and comp795(wire924, inA[24], inB[27]);
	and comp796(wire925, inA[24], inB[28]);
	and comp797(wire926, inA[24], inB[29]);
	and comp798(wire927, inA[24], inB[30]);
	and comp799(wire928, inA[24], inB[31]);
	and comp800(wire929, inA[25], inB[0]);
	and comp801(wire930, inA[25], inB[1]);
	and comp802(wire931, inA[25], inB[2]);
	and comp803(wire932, inA[25], inB[3]);
	and comp804(wire933, inA[25], inB[4]);
	and comp805(wire934, inA[25], inB[5]);
	and comp806(wire935, inA[25], inB[6]);
	and comp807(wire936, inA[25], inB[7]);
	and comp808(wire937, inA[25], inB[8]);
	and comp809(wire938, inA[25], inB[9]);
	and comp810(wire939, inA[25], inB[10]);
	and comp811(wire940, inA[25], inB[11]);
	and comp812(wire941, inA[25], inB[12]);
	and comp813(wire942, inA[25], inB[13]);
	and comp814(wire943, inA[25], inB[14]);
	and comp815(wire944, inA[25], inB[15]);
	and comp816(wire945, inA[25], inB[16]);
	and comp817(wire946, inA[25], inB[17]);
	and comp818(wire947, inA[25], inB[18]);
	and comp819(wire948, inA[25], inB[19]);
	and comp820(wire949, inA[25], inB[20]);
	and comp821(wire950, inA[25], inB[21]);
	and comp822(wire951, inA[25], inB[22]);
	and comp823(wire952, inA[25], inB[23]);
	and comp824(wire953, inA[25], inB[24]);
	and comp825(wire954, inA[25], inB[25]);
	and comp826(wire955, inA[25], inB[26]);
	and comp827(wire956, inA[25], inB[27]);
	and comp828(wire957, inA[25], inB[28]);
	and comp829(wire958, inA[25], inB[29]);
	and comp830(wire959, inA[25], inB[30]);
	and comp831(wire960, inA[25], inB[31]);
	and comp832(wire961, inA[26], inB[0]);
	and comp833(wire962, inA[26], inB[1]);
	and comp834(wire963, inA[26], inB[2]);
	and comp835(wire964, inA[26], inB[3]);
	and comp836(wire965, inA[26], inB[4]);
	and comp837(wire966, inA[26], inB[5]);
	and comp838(wire967, inA[26], inB[6]);
	and comp839(wire968, inA[26], inB[7]);
	and comp840(wire969, inA[26], inB[8]);
	and comp841(wire970, inA[26], inB[9]);
	and comp842(wire971, inA[26], inB[10]);
	and comp843(wire972, inA[26], inB[11]);
	and comp844(wire973, inA[26], inB[12]);
	and comp845(wire974, inA[26], inB[13]);
	and comp846(wire975, inA[26], inB[14]);
	and comp847(wire976, inA[26], inB[15]);
	and comp848(wire977, inA[26], inB[16]);
	and comp849(wire978, inA[26], inB[17]);
	and comp850(wire979, inA[26], inB[18]);
	and comp851(wire980, inA[26], inB[19]);
	and comp852(wire981, inA[26], inB[20]);
	and comp853(wire982, inA[26], inB[21]);
	and comp854(wire983, inA[26], inB[22]);
	and comp855(wire984, inA[26], inB[23]);
	and comp856(wire985, inA[26], inB[24]);
	and comp857(wire986, inA[26], inB[25]);
	and comp858(wire987, inA[26], inB[26]);
	and comp859(wire988, inA[26], inB[27]);
	and comp860(wire989, inA[26], inB[28]);
	and comp861(wire990, inA[26], inB[29]);
	and comp862(wire991, inA[26], inB[30]);
	and comp863(wire992, inA[26], inB[31]);
	and comp864(wire993, inA[27], inB[0]);
	and comp865(wire994, inA[27], inB[1]);
	and comp866(wire995, inA[27], inB[2]);
	and comp867(wire996, inA[27], inB[3]);
	and comp868(wire997, inA[27], inB[4]);
	and comp869(wire998, inA[27], inB[5]);
	and comp870(wire999, inA[27], inB[6]);
	and comp871(wire1000, inA[27], inB[7]);
	and comp872(wire1001, inA[27], inB[8]);
	and comp873(wire1002, inA[27], inB[9]);
	and comp874(wire1003, inA[27], inB[10]);
	and comp875(wire1004, inA[27], inB[11]);
	and comp876(wire1005, inA[27], inB[12]);
	and comp877(wire1006, inA[27], inB[13]);
	and comp878(wire1007, inA[27], inB[14]);
	and comp879(wire1008, inA[27], inB[15]);
	and comp880(wire1009, inA[27], inB[16]);
	and comp881(wire1010, inA[27], inB[17]);
	and comp882(wire1011, inA[27], inB[18]);
	and comp883(wire1012, inA[27], inB[19]);
	and comp884(wire1013, inA[27], inB[20]);
	and comp885(wire1014, inA[27], inB[21]);
	and comp886(wire1015, inA[27], inB[22]);
	and comp887(wire1016, inA[27], inB[23]);
	and comp888(wire1017, inA[27], inB[24]);
	and comp889(wire1018, inA[27], inB[25]);
	and comp890(wire1019, inA[27], inB[26]);
	and comp891(wire1020, inA[27], inB[27]);
	and comp892(wire1021, inA[27], inB[28]);
	and comp893(wire1022, inA[27], inB[29]);
	and comp894(wire1023, inA[27], inB[30]);
	and comp895(wire1024, inA[27], inB[31]);
	and comp896(wire1025, inA[28], inB[0]);
	and comp897(wire1026, inA[28], inB[1]);
	and comp898(wire1027, inA[28], inB[2]);
	and comp899(wire1028, inA[28], inB[3]);
	and comp900(wire1029, inA[28], inB[4]);
	and comp901(wire1030, inA[28], inB[5]);
	and comp902(wire1031, inA[28], inB[6]);
	and comp903(wire1032, inA[28], inB[7]);
	and comp904(wire1033, inA[28], inB[8]);
	and comp905(wire1034, inA[28], inB[9]);
	and comp906(wire1035, inA[28], inB[10]);
	and comp907(wire1036, inA[28], inB[11]);
	and comp908(wire1037, inA[28], inB[12]);
	and comp909(wire1038, inA[28], inB[13]);
	and comp910(wire1039, inA[28], inB[14]);
	and comp911(wire1040, inA[28], inB[15]);
	and comp912(wire1041, inA[28], inB[16]);
	and comp913(wire1042, inA[28], inB[17]);
	and comp914(wire1043, inA[28], inB[18]);
	and comp915(wire1044, inA[28], inB[19]);
	and comp916(wire1045, inA[28], inB[20]);
	and comp917(wire1046, inA[28], inB[21]);
	and comp918(wire1047, inA[28], inB[22]);
	and comp919(wire1048, inA[28], inB[23]);
	and comp920(wire1049, inA[28], inB[24]);
	and comp921(wire1050, inA[28], inB[25]);
	and comp922(wire1051, inA[28], inB[26]);
	and comp923(wire1052, inA[28], inB[27]);
	and comp924(wire1053, inA[28], inB[28]);
	and comp925(wire1054, inA[28], inB[29]);
	and comp926(wire1055, inA[28], inB[30]);
	and comp927(wire1056, inA[28], inB[31]);
	and comp928(wire1057, inA[29], inB[0]);
	and comp929(wire1058, inA[29], inB[1]);
	and comp930(wire1059, inA[29], inB[2]);
	and comp931(wire1060, inA[29], inB[3]);
	and comp932(wire1061, inA[29], inB[4]);
	and comp933(wire1062, inA[29], inB[5]);
	and comp934(wire1063, inA[29], inB[6]);
	and comp935(wire1064, inA[29], inB[7]);
	and comp936(wire1065, inA[29], inB[8]);
	and comp937(wire1066, inA[29], inB[9]);
	and comp938(wire1067, inA[29], inB[10]);
	and comp939(wire1068, inA[29], inB[11]);
	and comp940(wire1069, inA[29], inB[12]);
	and comp941(wire1070, inA[29], inB[13]);
	and comp942(wire1071, inA[29], inB[14]);
	and comp943(wire1072, inA[29], inB[15]);
	and comp944(wire1073, inA[29], inB[16]);
	and comp945(wire1074, inA[29], inB[17]);
	and comp946(wire1075, inA[29], inB[18]);
	and comp947(wire1076, inA[29], inB[19]);
	and comp948(wire1077, inA[29], inB[20]);
	and comp949(wire1078, inA[29], inB[21]);
	and comp950(wire1079, inA[29], inB[22]);
	and comp951(wire1080, inA[29], inB[23]);
	and comp952(wire1081, inA[29], inB[24]);
	and comp953(wire1082, inA[29], inB[25]);
	and comp954(wire1083, inA[29], inB[26]);
	and comp955(wire1084, inA[29], inB[27]);
	and comp956(wire1085, inA[29], inB[28]);
	and comp957(wire1086, inA[29], inB[29]);
	and comp958(wire1087, inA[29], inB[30]);
	and comp959(wire1088, inA[29], inB[31]);
	and comp960(wire1089, inA[30], inB[0]);
	and comp961(wire1090, inA[30], inB[1]);
	and comp962(wire1091, inA[30], inB[2]);
	and comp963(wire1092, inA[30], inB[3]);
	and comp964(wire1093, inA[30], inB[4]);
	and comp965(wire1094, inA[30], inB[5]);
	and comp966(wire1095, inA[30], inB[6]);
	and comp967(wire1096, inA[30], inB[7]);
	and comp968(wire1097, inA[30], inB[8]);
	and comp969(wire1098, inA[30], inB[9]);
	and comp970(wire1099, inA[30], inB[10]);
	and comp971(wire1100, inA[30], inB[11]);
	and comp972(wire1101, inA[30], inB[12]);
	and comp973(wire1102, inA[30], inB[13]);
	and comp974(wire1103, inA[30], inB[14]);
	and comp975(wire1104, inA[30], inB[15]);
	and comp976(wire1105, inA[30], inB[16]);
	and comp977(wire1106, inA[30], inB[17]);
	and comp978(wire1107, inA[30], inB[18]);
	and comp979(wire1108, inA[30], inB[19]);
	and comp980(wire1109, inA[30], inB[20]);
	and comp981(wire1110, inA[30], inB[21]);
	and comp982(wire1111, inA[30], inB[22]);
	and comp983(wire1112, inA[30], inB[23]);
	and comp984(wire1113, inA[30], inB[24]);
	and comp985(wire1114, inA[30], inB[25]);
	and comp986(wire1115, inA[30], inB[26]);
	and comp987(wire1116, inA[30], inB[27]);
	and comp988(wire1117, inA[30], inB[28]);
	and comp989(wire1118, inA[30], inB[29]);
	and comp990(wire1119, inA[30], inB[30]);
	and comp991(wire1120, inA[30], inB[31]);
	and comp992(wire1121, inA[31], inB[0]);
	and comp993(wire1122, inA[31], inB[1]);
	and comp994(wire1123, inA[31], inB[2]);
	and comp995(wire1124, inA[31], inB[3]);
	and comp996(wire1125, inA[31], inB[4]);
	and comp997(wire1126, inA[31], inB[5]);
	and comp998(wire1127, inA[31], inB[6]);
	and comp999(wire1128, inA[31], inB[7]);
	and comp1000(wire1129, inA[31], inB[8]);
	and comp1001(wire1130, inA[31], inB[9]);
	and comp1002(wire1131, inA[31], inB[10]);
	and comp1003(wire1132, inA[31], inB[11]);
	and comp1004(wire1133, inA[31], inB[12]);
	and comp1005(wire1134, inA[31], inB[13]);
	and comp1006(wire1135, inA[31], inB[14]);
	and comp1007(wire1136, inA[31], inB[15]);
	and comp1008(wire1137, inA[31], inB[16]);
	and comp1009(wire1138, inA[31], inB[17]);
	and comp1010(wire1139, inA[31], inB[18]);
	and comp1011(wire1140, inA[31], inB[19]);
	and comp1012(wire1141, inA[31], inB[20]);
	and comp1013(wire1142, inA[31], inB[21]);
	and comp1014(wire1143, inA[31], inB[22]);
	and comp1015(wire1144, inA[31], inB[23]);
	and comp1016(wire1145, inA[31], inB[24]);
	and comp1017(wire1146, inA[31], inB[25]);
	and comp1018(wire1147, inA[31], inB[26]);
	and comp1019(wire1148, inA[31], inB[27]);
	and comp1020(wire1149, inA[31], inB[28]);
	and comp1021(wire1150, inA[31], inB[29]);
	and comp1022(wire1151, inA[31], inB[30]);
	and comp1023(wire1152, inA[31], inB[31]);
	half_add comp1024(.out(wire1153), .cout(wire1154), .inA(wire157), .inB(wire188));
	full_add comp1025(.out(wire1155), .cout(wire1156), .inA(wire158), .inB(wire189), .cin(wire220));
	half_add comp1026(.out(wire1157), .cout(wire1158), .inA(wire251), .inB(wire282));
	full_add comp1027(.out(wire1159), .cout(wire1160), .inA(wire159), .inB(wire190), .cin(wire221));
	full_add comp1028(.out(wire1161), .cout(wire1162), .inA(wire252), .inB(wire283), .cin(wire314));
	half_add comp1029(.out(wire1163), .cout(wire1164), .inA(wire345), .inB(wire376));
	full_add comp1030(.out(wire1165), .cout(wire1166), .inA(wire160), .inB(wire191), .cin(wire222));
	full_add comp1031(.out(wire1167), .cout(wire1168), .inA(wire253), .inB(wire284), .cin(wire315));
	full_add comp1032(.out(wire1169), .cout(wire1170), .inA(wire346), .inB(wire377), .cin(wire408));
	half_add comp1033(.out(wire1171), .cout(wire1172), .inA(wire439), .inB(wire470));
	full_add comp1034(.out(wire1173), .cout(wire1174), .inA(wire192), .inB(wire223), .cin(wire254));
	full_add comp1035(.out(wire1175), .cout(wire1176), .inA(wire285), .inB(wire316), .cin(wire347));
	full_add comp1036(.out(wire1177), .cout(wire1178), .inA(wire378), .inB(wire409), .cin(wire440));
	half_add comp1037(.out(wire1179), .cout(wire1180), .inA(wire471), .inB(wire502));
	full_add comp1038(.out(wire1181), .cout(wire1182), .inA(wire224), .inB(wire255), .cin(wire286));
	full_add comp1039(.out(wire1183), .cout(wire1184), .inA(wire317), .inB(wire348), .cin(wire379));
	full_add comp1040(.out(wire1185), .cout(wire1186), .inA(wire410), .inB(wire441), .cin(wire472));
	full_add comp1041(.out(wire1187), .cout(wire1188), .inA(wire256), .inB(wire287), .cin(wire318));
	full_add comp1042(.out(wire1189), .cout(wire1190), .inA(wire349), .inB(wire380), .cin(wire411));
	full_add comp1043(.out(wire1191), .cout(wire1192), .inA(wire288), .inB(wire319), .cin(wire350));
	half_add comp1044(.out(wire1193), .cout(wire1194), .inA(wire148), .inB(wire179));
	full_add comp1045(.out(wire1195), .cout(wire1196), .inA(wire149), .inB(wire180), .cin(wire211));
	half_add comp1046(.out(wire1197), .cout(wire1198), .inA(wire242), .inB(wire273));
	full_add comp1047(.out(wire1199), .cout(wire1200), .inA(wire150), .inB(wire181), .cin(wire212));
	full_add comp1048(.out(wire1201), .cout(wire1202), .inA(wire243), .inB(wire274), .cin(wire305));
	half_add comp1049(.out(wire1203), .cout(wire1204), .inA(wire336), .inB(wire367));
	full_add comp1050(.out(wire1205), .cout(wire1206), .inA(wire151), .inB(wire182), .cin(wire213));
	full_add comp1051(.out(wire1207), .cout(wire1208), .inA(wire244), .inB(wire275), .cin(wire306));
	full_add comp1052(.out(wire1209), .cout(wire1210), .inA(wire337), .inB(wire368), .cin(wire399));
	half_add comp1053(.out(wire1211), .cout(wire1212), .inA(wire430), .inB(wire461));
	full_add comp1054(.out(wire1213), .cout(wire1214), .inA(wire152), .inB(wire183), .cin(wire214));
	full_add comp1055(.out(wire1215), .cout(wire1216), .inA(wire245), .inB(wire276), .cin(wire307));
	full_add comp1056(.out(wire1217), .cout(wire1218), .inA(wire338), .inB(wire369), .cin(wire400));
	full_add comp1057(.out(wire1219), .cout(wire1220), .inA(wire431), .inB(wire462), .cin(wire493));
	half_add comp1058(.out(wire1221), .cout(wire1222), .inA(wire524), .inB(wire555));
	full_add comp1059(.out(wire1223), .cout(wire1224), .inA(wire153), .inB(wire184), .cin(wire215));
	full_add comp1060(.out(wire1225), .cout(wire1226), .inA(wire246), .inB(wire277), .cin(wire308));
	full_add comp1061(.out(wire1227), .cout(wire1228), .inA(wire339), .inB(wire370), .cin(wire401));
	full_add comp1062(.out(wire1229), .cout(wire1230), .inA(wire432), .inB(wire463), .cin(wire494));
	full_add comp1063(.out(wire1231), .cout(wire1232), .inA(wire525), .inB(wire556), .cin(wire587));
	half_add comp1064(.out(wire1233), .cout(wire1234), .inA(wire618), .inB(wire649));
	full_add comp1065(.out(wire1235), .cout(wire1236), .inA(wire154), .inB(wire185), .cin(wire216));
	full_add comp1066(.out(wire1237), .cout(wire1238), .inA(wire247), .inB(wire278), .cin(wire309));
	full_add comp1067(.out(wire1239), .cout(wire1240), .inA(wire340), .inB(wire371), .cin(wire402));
	full_add comp1068(.out(wire1241), .cout(wire1242), .inA(wire433), .inB(wire464), .cin(wire495));
	full_add comp1069(.out(wire1243), .cout(wire1244), .inA(wire526), .inB(wire557), .cin(wire588));
	full_add comp1070(.out(wire1245), .cout(wire1246), .inA(wire619), .inB(wire650), .cin(wire681));
	half_add comp1071(.out(wire1247), .cout(wire1248), .inA(wire712), .inB(wire743));
	full_add comp1072(.out(wire1249), .cout(wire1250), .inA(wire155), .inB(wire186), .cin(wire217));
	full_add comp1073(.out(wire1251), .cout(wire1252), .inA(wire248), .inB(wire279), .cin(wire310));
	full_add comp1074(.out(wire1253), .cout(wire1254), .inA(wire341), .inB(wire372), .cin(wire403));
	full_add comp1075(.out(wire1255), .cout(wire1256), .inA(wire434), .inB(wire465), .cin(wire496));
	full_add comp1076(.out(wire1257), .cout(wire1258), .inA(wire527), .inB(wire558), .cin(wire589));
	full_add comp1077(.out(wire1259), .cout(wire1260), .inA(wire620), .inB(wire651), .cin(wire682));
	full_add comp1078(.out(wire1261), .cout(wire1262), .inA(wire713), .inB(wire744), .cin(wire775));
	half_add comp1079(.out(wire1263), .cout(wire1264), .inA(wire806), .inB(wire837));
	full_add comp1080(.out(wire1265), .cout(wire1266), .inA(wire156), .inB(wire187), .cin(wire218));
	full_add comp1081(.out(wire1267), .cout(wire1268), .inA(wire249), .inB(wire280), .cin(wire311));
	full_add comp1082(.out(wire1269), .cout(wire1270), .inA(wire342), .inB(wire373), .cin(wire404));
	full_add comp1083(.out(wire1271), .cout(wire1272), .inA(wire435), .inB(wire466), .cin(wire497));
	full_add comp1084(.out(wire1273), .cout(wire1274), .inA(wire528), .inB(wire559), .cin(wire590));
	full_add comp1085(.out(wire1275), .cout(wire1276), .inA(wire621), .inB(wire652), .cin(wire683));
	full_add comp1086(.out(wire1277), .cout(wire1278), .inA(wire714), .inB(wire745), .cin(wire776));
	full_add comp1087(.out(wire1279), .cout(wire1280), .inA(wire807), .inB(wire838), .cin(wire869));
	half_add comp1088(.out(wire1281), .cout(wire1282), .inA(wire900), .inB(wire931));
	full_add comp1089(.out(wire1283), .cout(wire1284), .inA(wire219), .inB(wire250), .cin(wire281));
	full_add comp1090(.out(wire1285), .cout(wire1286), .inA(wire312), .inB(wire343), .cin(wire374));
	full_add comp1091(.out(wire1287), .cout(wire1288), .inA(wire405), .inB(wire436), .cin(wire467));
	full_add comp1092(.out(wire1289), .cout(wire1290), .inA(wire498), .inB(wire529), .cin(wire560));
	full_add comp1093(.out(wire1291), .cout(wire1292), .inA(wire591), .inB(wire622), .cin(wire653));
	full_add comp1094(.out(wire1293), .cout(wire1294), .inA(wire684), .inB(wire715), .cin(wire746));
	full_add comp1095(.out(wire1295), .cout(wire1296), .inA(wire777), .inB(wire808), .cin(wire839));
	full_add comp1096(.out(wire1297), .cout(wire1298), .inA(wire870), .inB(wire901), .cin(wire932));
	full_add comp1097(.out(wire1299), .cout(wire1300), .inA(wire963), .inB(wire994), .cin(wire1025));
	full_add comp1098(.out(wire1301), .cout(wire1302), .inA(wire313), .inB(wire344), .cin(wire375));
	full_add comp1099(.out(wire1303), .cout(wire1304), .inA(wire406), .inB(wire437), .cin(wire468));
	full_add comp1100(.out(wire1305), .cout(wire1306), .inA(wire499), .inB(wire530), .cin(wire561));
	full_add comp1101(.out(wire1307), .cout(wire1308), .inA(wire592), .inB(wire623), .cin(wire654));
	full_add comp1102(.out(wire1309), .cout(wire1310), .inA(wire685), .inB(wire716), .cin(wire747));
	full_add comp1103(.out(wire1311), .cout(wire1312), .inA(wire778), .inB(wire809), .cin(wire840));
	full_add comp1104(.out(wire1313), .cout(wire1314), .inA(wire871), .inB(wire902), .cin(wire933));
	full_add comp1105(.out(wire1315), .cout(wire1316), .inA(wire964), .inB(wire995), .cin(wire1026));
	full_add comp1106(.out(wire1317), .cout(wire1318), .inA(wire1057), .inB(wire1154), .cin(wire1155));
	full_add comp1107(.out(wire1319), .cout(wire1320), .inA(wire407), .inB(wire438), .cin(wire469));
	full_add comp1108(.out(wire1321), .cout(wire1322), .inA(wire500), .inB(wire531), .cin(wire562));
	full_add comp1109(.out(wire1323), .cout(wire1324), .inA(wire593), .inB(wire624), .cin(wire655));
	full_add comp1110(.out(wire1325), .cout(wire1326), .inA(wire686), .inB(wire717), .cin(wire748));
	full_add comp1111(.out(wire1327), .cout(wire1328), .inA(wire779), .inB(wire810), .cin(wire841));
	full_add comp1112(.out(wire1329), .cout(wire1330), .inA(wire872), .inB(wire903), .cin(wire934));
	full_add comp1113(.out(wire1331), .cout(wire1332), .inA(wire965), .inB(wire996), .cin(wire1027));
	full_add comp1114(.out(wire1333), .cout(wire1334), .inA(wire1058), .inB(wire1089), .cin(wire1156));
	full_add comp1115(.out(wire1335), .cout(wire1336), .inA(wire1158), .inB(wire1159), .cin(wire1161));
	full_add comp1116(.out(wire1337), .cout(wire1338), .inA(wire501), .inB(wire532), .cin(wire563));
	full_add comp1117(.out(wire1339), .cout(wire1340), .inA(wire594), .inB(wire625), .cin(wire656));
	full_add comp1118(.out(wire1341), .cout(wire1342), .inA(wire687), .inB(wire718), .cin(wire749));
	full_add comp1119(.out(wire1343), .cout(wire1344), .inA(wire780), .inB(wire811), .cin(wire842));
	full_add comp1120(.out(wire1345), .cout(wire1346), .inA(wire873), .inB(wire904), .cin(wire935));
	full_add comp1121(.out(wire1347), .cout(wire1348), .inA(wire966), .inB(wire997), .cin(wire1028));
	full_add comp1122(.out(wire1349), .cout(wire1350), .inA(wire1059), .inB(wire1090), .cin(wire1121));
	full_add comp1123(.out(wire1351), .cout(wire1352), .inA(wire1160), .inB(wire1162), .cin(wire1164));
	full_add comp1124(.out(wire1353), .cout(wire1354), .inA(wire1165), .inB(wire1167), .cin(wire1169));
	full_add comp1125(.out(wire1355), .cout(wire1356), .inA(wire533), .inB(wire564), .cin(wire595));
	full_add comp1126(.out(wire1357), .cout(wire1358), .inA(wire626), .inB(wire657), .cin(wire688));
	full_add comp1127(.out(wire1359), .cout(wire1360), .inA(wire719), .inB(wire750), .cin(wire781));
	full_add comp1128(.out(wire1361), .cout(wire1362), .inA(wire812), .inB(wire843), .cin(wire874));
	full_add comp1129(.out(wire1363), .cout(wire1364), .inA(wire905), .inB(wire936), .cin(wire967));
	full_add comp1130(.out(wire1365), .cout(wire1366), .inA(wire998), .inB(wire1029), .cin(wire1060));
	full_add comp1131(.out(wire1367), .cout(wire1368), .inA(wire1091), .inB(wire1122), .cin(wire1166));
	full_add comp1132(.out(wire1369), .cout(wire1370), .inA(wire1168), .inB(wire1170), .cin(wire1172));
	full_add comp1133(.out(wire1371), .cout(wire1372), .inA(wire1173), .inB(wire1175), .cin(wire1177));
	full_add comp1134(.out(wire1373), .cout(wire1374), .inA(wire503), .inB(wire534), .cin(wire565));
	full_add comp1135(.out(wire1375), .cout(wire1376), .inA(wire596), .inB(wire627), .cin(wire658));
	full_add comp1136(.out(wire1377), .cout(wire1378), .inA(wire689), .inB(wire720), .cin(wire751));
	full_add comp1137(.out(wire1379), .cout(wire1380), .inA(wire782), .inB(wire813), .cin(wire844));
	full_add comp1138(.out(wire1381), .cout(wire1382), .inA(wire875), .inB(wire906), .cin(wire937));
	full_add comp1139(.out(wire1383), .cout(wire1384), .inA(wire968), .inB(wire999), .cin(wire1030));
	full_add comp1140(.out(wire1385), .cout(wire1386), .inA(wire1061), .inB(wire1092), .cin(wire1123));
	full_add comp1141(.out(wire1387), .cout(wire1388), .inA(wire1174), .inB(wire1176), .cin(wire1178));
	full_add comp1142(.out(wire1389), .cout(wire1390), .inA(wire1180), .inB(wire1181), .cin(wire1183));
	full_add comp1143(.out(wire1391), .cout(wire1392), .inA(wire442), .inB(wire473), .cin(wire504));
	full_add comp1144(.out(wire1393), .cout(wire1394), .inA(wire535), .inB(wire566), .cin(wire597));
	full_add comp1145(.out(wire1395), .cout(wire1396), .inA(wire628), .inB(wire659), .cin(wire690));
	full_add comp1146(.out(wire1397), .cout(wire1398), .inA(wire721), .inB(wire752), .cin(wire783));
	full_add comp1147(.out(wire1399), .cout(wire1400), .inA(wire814), .inB(wire845), .cin(wire876));
	full_add comp1148(.out(wire1401), .cout(wire1402), .inA(wire907), .inB(wire938), .cin(wire969));
	full_add comp1149(.out(wire1403), .cout(wire1404), .inA(wire1000), .inB(wire1031), .cin(wire1062));
	full_add comp1150(.out(wire1405), .cout(wire1406), .inA(wire1093), .inB(wire1124), .cin(wire1182));
	full_add comp1151(.out(wire1407), .cout(wire1408), .inA(wire1184), .inB(wire1186), .cin(wire1187));
	full_add comp1152(.out(wire1409), .cout(wire1410), .inA(wire381), .inB(wire412), .cin(wire443));
	full_add comp1153(.out(wire1411), .cout(wire1412), .inA(wire474), .inB(wire505), .cin(wire536));
	full_add comp1154(.out(wire1413), .cout(wire1414), .inA(wire567), .inB(wire598), .cin(wire629));
	full_add comp1155(.out(wire1415), .cout(wire1416), .inA(wire660), .inB(wire691), .cin(wire722));
	full_add comp1156(.out(wire1417), .cout(wire1418), .inA(wire753), .inB(wire784), .cin(wire815));
	full_add comp1157(.out(wire1419), .cout(wire1420), .inA(wire846), .inB(wire877), .cin(wire908));
	full_add comp1158(.out(wire1421), .cout(wire1422), .inA(wire939), .inB(wire970), .cin(wire1001));
	full_add comp1159(.out(wire1423), .cout(wire1424), .inA(wire1032), .inB(wire1063), .cin(wire1094));
	full_add comp1160(.out(wire1425), .cout(wire1426), .inA(wire1125), .inB(wire1188), .cin(wire1190));
	full_add comp1161(.out(wire1427), .cout(wire1428), .inA(wire320), .inB(wire351), .cin(wire382));
	full_add comp1162(.out(wire1429), .cout(wire1430), .inA(wire413), .inB(wire444), .cin(wire475));
	full_add comp1163(.out(wire1431), .cout(wire1432), .inA(wire506), .inB(wire537), .cin(wire568));
	full_add comp1164(.out(wire1433), .cout(wire1434), .inA(wire599), .inB(wire630), .cin(wire661));
	full_add comp1165(.out(wire1435), .cout(wire1436), .inA(wire692), .inB(wire723), .cin(wire754));
	full_add comp1166(.out(wire1437), .cout(wire1438), .inA(wire785), .inB(wire816), .cin(wire847));
	full_add comp1167(.out(wire1439), .cout(wire1440), .inA(wire878), .inB(wire909), .cin(wire940));
	full_add comp1168(.out(wire1441), .cout(wire1442), .inA(wire971), .inB(wire1002), .cin(wire1033));
	full_add comp1169(.out(wire1443), .cout(wire1444), .inA(wire1064), .inB(wire1095), .cin(wire1126));
	full_add comp1170(.out(wire1445), .cout(wire1446), .inA(wire352), .inB(wire383), .cin(wire414));
	full_add comp1171(.out(wire1447), .cout(wire1448), .inA(wire445), .inB(wire476), .cin(wire507));
	full_add comp1172(.out(wire1449), .cout(wire1450), .inA(wire538), .inB(wire569), .cin(wire600));
	full_add comp1173(.out(wire1451), .cout(wire1452), .inA(wire631), .inB(wire662), .cin(wire693));
	full_add comp1174(.out(wire1453), .cout(wire1454), .inA(wire724), .inB(wire755), .cin(wire786));
	full_add comp1175(.out(wire1455), .cout(wire1456), .inA(wire817), .inB(wire848), .cin(wire879));
	full_add comp1176(.out(wire1457), .cout(wire1458), .inA(wire910), .inB(wire941), .cin(wire972));
	full_add comp1177(.out(wire1459), .cout(wire1460), .inA(wire1003), .inB(wire1034), .cin(wire1065));
	full_add comp1178(.out(wire1461), .cout(wire1462), .inA(wire384), .inB(wire415), .cin(wire446));
	full_add comp1179(.out(wire1463), .cout(wire1464), .inA(wire477), .inB(wire508), .cin(wire539));
	full_add comp1180(.out(wire1465), .cout(wire1466), .inA(wire570), .inB(wire601), .cin(wire632));
	full_add comp1181(.out(wire1467), .cout(wire1468), .inA(wire663), .inB(wire694), .cin(wire725));
	full_add comp1182(.out(wire1469), .cout(wire1470), .inA(wire756), .inB(wire787), .cin(wire818));
	full_add comp1183(.out(wire1471), .cout(wire1472), .inA(wire849), .inB(wire880), .cin(wire911));
	full_add comp1184(.out(wire1473), .cout(wire1474), .inA(wire942), .inB(wire973), .cin(wire1004));
	full_add comp1185(.out(wire1475), .cout(wire1476), .inA(wire416), .inB(wire447), .cin(wire478));
	full_add comp1186(.out(wire1477), .cout(wire1478), .inA(wire509), .inB(wire540), .cin(wire571));
	full_add comp1187(.out(wire1479), .cout(wire1480), .inA(wire602), .inB(wire633), .cin(wire664));
	full_add comp1188(.out(wire1481), .cout(wire1482), .inA(wire695), .inB(wire726), .cin(wire757));
	full_add comp1189(.out(wire1483), .cout(wire1484), .inA(wire788), .inB(wire819), .cin(wire850));
	full_add comp1190(.out(wire1485), .cout(wire1486), .inA(wire881), .inB(wire912), .cin(wire943));
	full_add comp1191(.out(wire1487), .cout(wire1488), .inA(wire448), .inB(wire479), .cin(wire510));
	full_add comp1192(.out(wire1489), .cout(wire1490), .inA(wire541), .inB(wire572), .cin(wire603));
	full_add comp1193(.out(wire1491), .cout(wire1492), .inA(wire634), .inB(wire665), .cin(wire696));
	full_add comp1194(.out(wire1493), .cout(wire1494), .inA(wire727), .inB(wire758), .cin(wire789));
	full_add comp1195(.out(wire1495), .cout(wire1496), .inA(wire820), .inB(wire851), .cin(wire882));
	full_add comp1196(.out(wire1497), .cout(wire1498), .inA(wire480), .inB(wire511), .cin(wire542));
	full_add comp1197(.out(wire1499), .cout(wire1500), .inA(wire573), .inB(wire604), .cin(wire635));
	full_add comp1198(.out(wire1501), .cout(wire1502), .inA(wire666), .inB(wire697), .cin(wire728));
	full_add comp1199(.out(wire1503), .cout(wire1504), .inA(wire759), .inB(wire790), .cin(wire821));
	full_add comp1200(.out(wire1505), .cout(wire1506), .inA(wire512), .inB(wire543), .cin(wire574));
	full_add comp1201(.out(wire1507), .cout(wire1508), .inA(wire605), .inB(wire636), .cin(wire667));
	full_add comp1202(.out(wire1509), .cout(wire1510), .inA(wire698), .inB(wire729), .cin(wire760));
	full_add comp1203(.out(wire1511), .cout(wire1512), .inA(wire544), .inB(wire575), .cin(wire606));
	full_add comp1204(.out(wire1513), .cout(wire1514), .inA(wire637), .inB(wire668), .cin(wire699));
	full_add comp1205(.out(wire1515), .cout(wire1516), .inA(wire576), .inB(wire607), .cin(wire638));
	half_add comp1206(.out(wire1517), .cout(wire1518), .inA(wire142), .inB(wire173));
	full_add comp1207(.out(wire1519), .cout(wire1520), .inA(wire143), .inB(wire174), .cin(wire205));
	half_add comp1208(.out(wire1521), .cout(wire1522), .inA(wire236), .inB(wire267));
	full_add comp1209(.out(wire1523), .cout(wire1524), .inA(wire144), .inB(wire175), .cin(wire206));
	full_add comp1210(.out(wire1525), .cout(wire1526), .inA(wire237), .inB(wire268), .cin(wire299));
	half_add comp1211(.out(wire1527), .cout(wire1528), .inA(wire330), .inB(wire361));
	full_add comp1212(.out(wire1529), .cout(wire1530), .inA(wire145), .inB(wire176), .cin(wire207));
	full_add comp1213(.out(wire1531), .cout(wire1532), .inA(wire238), .inB(wire269), .cin(wire300));
	full_add comp1214(.out(wire1533), .cout(wire1534), .inA(wire331), .inB(wire362), .cin(wire393));
	half_add comp1215(.out(wire1535), .cout(wire1536), .inA(wire424), .inB(wire455));
	full_add comp1216(.out(wire1537), .cout(wire1538), .inA(wire146), .inB(wire177), .cin(wire208));
	full_add comp1217(.out(wire1539), .cout(wire1540), .inA(wire239), .inB(wire270), .cin(wire301));
	full_add comp1218(.out(wire1541), .cout(wire1542), .inA(wire332), .inB(wire363), .cin(wire394));
	full_add comp1219(.out(wire1543), .cout(wire1544), .inA(wire425), .inB(wire456), .cin(wire487));
	half_add comp1220(.out(wire1545), .cout(wire1546), .inA(wire518), .inB(wire549));
	full_add comp1221(.out(wire1547), .cout(wire1548), .inA(wire147), .inB(wire178), .cin(wire209));
	full_add comp1222(.out(wire1549), .cout(wire1550), .inA(wire240), .inB(wire271), .cin(wire302));
	full_add comp1223(.out(wire1551), .cout(wire1552), .inA(wire333), .inB(wire364), .cin(wire395));
	full_add comp1224(.out(wire1553), .cout(wire1554), .inA(wire426), .inB(wire457), .cin(wire488));
	full_add comp1225(.out(wire1555), .cout(wire1556), .inA(wire519), .inB(wire550), .cin(wire581));
	half_add comp1226(.out(wire1557), .cout(wire1558), .inA(wire612), .inB(wire643));
	full_add comp1227(.out(wire1559), .cout(wire1560), .inA(wire210), .inB(wire241), .cin(wire272));
	full_add comp1228(.out(wire1561), .cout(wire1562), .inA(wire303), .inB(wire334), .cin(wire365));
	full_add comp1229(.out(wire1563), .cout(wire1564), .inA(wire396), .inB(wire427), .cin(wire458));
	full_add comp1230(.out(wire1565), .cout(wire1566), .inA(wire489), .inB(wire520), .cin(wire551));
	full_add comp1231(.out(wire1567), .cout(wire1568), .inA(wire582), .inB(wire613), .cin(wire644));
	full_add comp1232(.out(wire1569), .cout(wire1570), .inA(wire675), .inB(wire706), .cin(wire737));
	full_add comp1233(.out(wire1571), .cout(wire1572), .inA(wire304), .inB(wire335), .cin(wire366));
	full_add comp1234(.out(wire1573), .cout(wire1574), .inA(wire397), .inB(wire428), .cin(wire459));
	full_add comp1235(.out(wire1575), .cout(wire1576), .inA(wire490), .inB(wire521), .cin(wire552));
	full_add comp1236(.out(wire1577), .cout(wire1578), .inA(wire583), .inB(wire614), .cin(wire645));
	full_add comp1237(.out(wire1579), .cout(wire1580), .inA(wire676), .inB(wire707), .cin(wire738));
	full_add comp1238(.out(wire1581), .cout(wire1582), .inA(wire769), .inB(wire1194), .cin(wire1195));
	full_add comp1239(.out(wire1583), .cout(wire1584), .inA(wire398), .inB(wire429), .cin(wire460));
	full_add comp1240(.out(wire1585), .cout(wire1586), .inA(wire491), .inB(wire522), .cin(wire553));
	full_add comp1241(.out(wire1587), .cout(wire1588), .inA(wire584), .inB(wire615), .cin(wire646));
	full_add comp1242(.out(wire1589), .cout(wire1590), .inA(wire677), .inB(wire708), .cin(wire739));
	full_add comp1243(.out(wire1591), .cout(wire1592), .inA(wire770), .inB(wire801), .cin(wire1196));
	full_add comp1244(.out(wire1593), .cout(wire1594), .inA(wire1198), .inB(wire1199), .cin(wire1201));
	full_add comp1245(.out(wire1595), .cout(wire1596), .inA(wire492), .inB(wire523), .cin(wire554));
	full_add comp1246(.out(wire1597), .cout(wire1598), .inA(wire585), .inB(wire616), .cin(wire647));
	full_add comp1247(.out(wire1599), .cout(wire1600), .inA(wire678), .inB(wire709), .cin(wire740));
	full_add comp1248(.out(wire1601), .cout(wire1602), .inA(wire771), .inB(wire802), .cin(wire833));
	full_add comp1249(.out(wire1603), .cout(wire1604), .inA(wire1200), .inB(wire1202), .cin(wire1204));
	full_add comp1250(.out(wire1605), .cout(wire1606), .inA(wire1205), .inB(wire1207), .cin(wire1209));
	full_add comp1251(.out(wire1607), .cout(wire1608), .inA(wire586), .inB(wire617), .cin(wire648));
	full_add comp1252(.out(wire1609), .cout(wire1610), .inA(wire679), .inB(wire710), .cin(wire741));
	full_add comp1253(.out(wire1611), .cout(wire1612), .inA(wire772), .inB(wire803), .cin(wire834));
	full_add comp1254(.out(wire1613), .cout(wire1614), .inA(wire865), .inB(wire1206), .cin(wire1208));
	full_add comp1255(.out(wire1615), .cout(wire1616), .inA(wire1210), .inB(wire1212), .cin(wire1213));
	full_add comp1256(.out(wire1617), .cout(wire1618), .inA(wire1215), .inB(wire1217), .cin(wire1219));
	full_add comp1257(.out(wire1619), .cout(wire1620), .inA(wire680), .inB(wire711), .cin(wire742));
	full_add comp1258(.out(wire1621), .cout(wire1622), .inA(wire773), .inB(wire804), .cin(wire835));
	full_add comp1259(.out(wire1623), .cout(wire1624), .inA(wire866), .inB(wire897), .cin(wire1214));
	full_add comp1260(.out(wire1625), .cout(wire1626), .inA(wire1216), .inB(wire1218), .cin(wire1220));
	full_add comp1261(.out(wire1627), .cout(wire1628), .inA(wire1222), .inB(wire1223), .cin(wire1225));
	full_add comp1262(.out(wire1629), .cout(wire1630), .inA(wire1227), .inB(wire1229), .cin(wire1231));
	full_add comp1263(.out(wire1631), .cout(wire1632), .inA(wire774), .inB(wire805), .cin(wire836));
	full_add comp1264(.out(wire1633), .cout(wire1634), .inA(wire867), .inB(wire898), .cin(wire929));
	full_add comp1265(.out(wire1635), .cout(wire1636), .inA(wire1224), .inB(wire1226), .cin(wire1228));
	full_add comp1266(.out(wire1637), .cout(wire1638), .inA(wire1230), .inB(wire1232), .cin(wire1234));
	full_add comp1267(.out(wire1639), .cout(wire1640), .inA(wire1235), .inB(wire1237), .cin(wire1239));
	full_add comp1268(.out(wire1641), .cout(wire1642), .inA(wire1241), .inB(wire1243), .cin(wire1245));
	full_add comp1269(.out(wire1643), .cout(wire1644), .inA(wire868), .inB(wire899), .cin(wire930));
	full_add comp1270(.out(wire1645), .cout(wire1646), .inA(wire961), .inB(wire1236), .cin(wire1238));
	full_add comp1271(.out(wire1647), .cout(wire1648), .inA(wire1240), .inB(wire1242), .cin(wire1244));
	full_add comp1272(.out(wire1649), .cout(wire1650), .inA(wire1246), .inB(wire1248), .cin(wire1249));
	full_add comp1273(.out(wire1651), .cout(wire1652), .inA(wire1251), .inB(wire1253), .cin(wire1255));
	full_add comp1274(.out(wire1653), .cout(wire1654), .inA(wire1257), .inB(wire1259), .cin(wire1261));
	full_add comp1275(.out(wire1655), .cout(wire1656), .inA(wire962), .inB(wire993), .cin(wire1250));
	full_add comp1276(.out(wire1657), .cout(wire1658), .inA(wire1252), .inB(wire1254), .cin(wire1256));
	full_add comp1277(.out(wire1659), .cout(wire1660), .inA(wire1258), .inB(wire1260), .cin(wire1262));
	full_add comp1278(.out(wire1661), .cout(wire1662), .inA(wire1264), .inB(wire1265), .cin(wire1267));
	full_add comp1279(.out(wire1663), .cout(wire1664), .inA(wire1269), .inB(wire1271), .cin(wire1273));
	full_add comp1280(.out(wire1665), .cout(wire1666), .inA(wire1275), .inB(wire1277), .cin(wire1279));
	full_add comp1281(.out(wire1667), .cout(wire1668), .inA(wire1153), .inB(wire1266), .cin(wire1268));
	full_add comp1282(.out(wire1669), .cout(wire1670), .inA(wire1270), .inB(wire1272), .cin(wire1274));
	full_add comp1283(.out(wire1671), .cout(wire1672), .inA(wire1276), .inB(wire1278), .cin(wire1280));
	full_add comp1284(.out(wire1673), .cout(wire1674), .inA(wire1282), .inB(wire1283), .cin(wire1285));
	full_add comp1285(.out(wire1675), .cout(wire1676), .inA(wire1287), .inB(wire1289), .cin(wire1291));
	full_add comp1286(.out(wire1677), .cout(wire1678), .inA(wire1293), .inB(wire1295), .cin(wire1297));
	full_add comp1287(.out(wire1679), .cout(wire1680), .inA(wire1157), .inB(wire1284), .cin(wire1286));
	full_add comp1288(.out(wire1681), .cout(wire1682), .inA(wire1288), .inB(wire1290), .cin(wire1292));
	full_add comp1289(.out(wire1683), .cout(wire1684), .inA(wire1294), .inB(wire1296), .cin(wire1298));
	full_add comp1290(.out(wire1685), .cout(wire1686), .inA(wire1300), .inB(wire1301), .cin(wire1303));
	full_add comp1291(.out(wire1687), .cout(wire1688), .inA(wire1305), .inB(wire1307), .cin(wire1309));
	full_add comp1292(.out(wire1689), .cout(wire1690), .inA(wire1311), .inB(wire1313), .cin(wire1315));
	full_add comp1293(.out(wire1691), .cout(wire1692), .inA(wire1163), .inB(wire1302), .cin(wire1304));
	full_add comp1294(.out(wire1693), .cout(wire1694), .inA(wire1306), .inB(wire1308), .cin(wire1310));
	full_add comp1295(.out(wire1695), .cout(wire1696), .inA(wire1312), .inB(wire1314), .cin(wire1316));
	full_add comp1296(.out(wire1697), .cout(wire1698), .inA(wire1318), .inB(wire1319), .cin(wire1321));
	full_add comp1297(.out(wire1699), .cout(wire1700), .inA(wire1323), .inB(wire1325), .cin(wire1327));
	full_add comp1298(.out(wire1701), .cout(wire1702), .inA(wire1329), .inB(wire1331), .cin(wire1333));
	full_add comp1299(.out(wire1703), .cout(wire1704), .inA(wire1171), .inB(wire1320), .cin(wire1322));
	full_add comp1300(.out(wire1705), .cout(wire1706), .inA(wire1324), .inB(wire1326), .cin(wire1328));
	full_add comp1301(.out(wire1707), .cout(wire1708), .inA(wire1330), .inB(wire1332), .cin(wire1334));
	full_add comp1302(.out(wire1709), .cout(wire1710), .inA(wire1336), .inB(wire1337), .cin(wire1339));
	full_add comp1303(.out(wire1711), .cout(wire1712), .inA(wire1341), .inB(wire1343), .cin(wire1345));
	full_add comp1304(.out(wire1713), .cout(wire1714), .inA(wire1347), .inB(wire1349), .cin(wire1351));
	full_add comp1305(.out(wire1715), .cout(wire1716), .inA(wire1179), .inB(wire1338), .cin(wire1340));
	full_add comp1306(.out(wire1717), .cout(wire1718), .inA(wire1342), .inB(wire1344), .cin(wire1346));
	full_add comp1307(.out(wire1719), .cout(wire1720), .inA(wire1348), .inB(wire1350), .cin(wire1352));
	full_add comp1308(.out(wire1721), .cout(wire1722), .inA(wire1354), .inB(wire1355), .cin(wire1357));
	full_add comp1309(.out(wire1723), .cout(wire1724), .inA(wire1359), .inB(wire1361), .cin(wire1363));
	full_add comp1310(.out(wire1725), .cout(wire1726), .inA(wire1365), .inB(wire1367), .cin(wire1369));
	full_add comp1311(.out(wire1727), .cout(wire1728), .inA(wire1185), .inB(wire1356), .cin(wire1358));
	full_add comp1312(.out(wire1729), .cout(wire1730), .inA(wire1360), .inB(wire1362), .cin(wire1364));
	full_add comp1313(.out(wire1731), .cout(wire1732), .inA(wire1366), .inB(wire1368), .cin(wire1370));
	full_add comp1314(.out(wire1733), .cout(wire1734), .inA(wire1372), .inB(wire1373), .cin(wire1375));
	full_add comp1315(.out(wire1735), .cout(wire1736), .inA(wire1377), .inB(wire1379), .cin(wire1381));
	full_add comp1316(.out(wire1737), .cout(wire1738), .inA(wire1383), .inB(wire1385), .cin(wire1387));
	full_add comp1317(.out(wire1739), .cout(wire1740), .inA(wire1189), .inB(wire1374), .cin(wire1376));
	full_add comp1318(.out(wire1741), .cout(wire1742), .inA(wire1378), .inB(wire1380), .cin(wire1382));
	full_add comp1319(.out(wire1743), .cout(wire1744), .inA(wire1384), .inB(wire1386), .cin(wire1388));
	full_add comp1320(.out(wire1745), .cout(wire1746), .inA(wire1390), .inB(wire1391), .cin(wire1393));
	full_add comp1321(.out(wire1747), .cout(wire1748), .inA(wire1395), .inB(wire1397), .cin(wire1399));
	full_add comp1322(.out(wire1749), .cout(wire1750), .inA(wire1401), .inB(wire1403), .cin(wire1405));
	full_add comp1323(.out(wire1751), .cout(wire1752), .inA(wire1191), .inB(wire1392), .cin(wire1394));
	full_add comp1324(.out(wire1753), .cout(wire1754), .inA(wire1396), .inB(wire1398), .cin(wire1400));
	full_add comp1325(.out(wire1755), .cout(wire1756), .inA(wire1402), .inB(wire1404), .cin(wire1406));
	full_add comp1326(.out(wire1757), .cout(wire1758), .inA(wire1408), .inB(wire1409), .cin(wire1411));
	full_add comp1327(.out(wire1759), .cout(wire1760), .inA(wire1413), .inB(wire1415), .cin(wire1417));
	full_add comp1328(.out(wire1761), .cout(wire1762), .inA(wire1419), .inB(wire1421), .cin(wire1423));
	full_add comp1329(.out(wire1763), .cout(wire1764), .inA(wire1192), .inB(wire1410), .cin(wire1412));
	full_add comp1330(.out(wire1765), .cout(wire1766), .inA(wire1414), .inB(wire1416), .cin(wire1418));
	full_add comp1331(.out(wire1767), .cout(wire1768), .inA(wire1420), .inB(wire1422), .cin(wire1424));
	full_add comp1332(.out(wire1769), .cout(wire1770), .inA(wire1426), .inB(wire1427), .cin(wire1429));
	full_add comp1333(.out(wire1771), .cout(wire1772), .inA(wire1431), .inB(wire1433), .cin(wire1435));
	full_add comp1334(.out(wire1773), .cout(wire1774), .inA(wire1437), .inB(wire1439), .cin(wire1441));
	full_add comp1335(.out(wire1775), .cout(wire1776), .inA(wire1096), .inB(wire1127), .cin(wire1428));
	full_add comp1336(.out(wire1777), .cout(wire1778), .inA(wire1430), .inB(wire1432), .cin(wire1434));
	full_add comp1337(.out(wire1779), .cout(wire1780), .inA(wire1436), .inB(wire1438), .cin(wire1440));
	full_add comp1338(.out(wire1781), .cout(wire1782), .inA(wire1442), .inB(wire1444), .cin(wire1445));
	full_add comp1339(.out(wire1783), .cout(wire1784), .inA(wire1447), .inB(wire1449), .cin(wire1451));
	full_add comp1340(.out(wire1785), .cout(wire1786), .inA(wire1453), .inB(wire1455), .cin(wire1457));
	full_add comp1341(.out(wire1787), .cout(wire1788), .inA(wire1035), .inB(wire1066), .cin(wire1097));
	full_add comp1342(.out(wire1789), .cout(wire1790), .inA(wire1128), .inB(wire1446), .cin(wire1448));
	full_add comp1343(.out(wire1791), .cout(wire1792), .inA(wire1450), .inB(wire1452), .cin(wire1454));
	full_add comp1344(.out(wire1793), .cout(wire1794), .inA(wire1456), .inB(wire1458), .cin(wire1460));
	full_add comp1345(.out(wire1795), .cout(wire1796), .inA(wire1461), .inB(wire1463), .cin(wire1465));
	full_add comp1346(.out(wire1797), .cout(wire1798), .inA(wire1467), .inB(wire1469), .cin(wire1471));
	full_add comp1347(.out(wire1799), .cout(wire1800), .inA(wire974), .inB(wire1005), .cin(wire1036));
	full_add comp1348(.out(wire1801), .cout(wire1802), .inA(wire1067), .inB(wire1098), .cin(wire1129));
	full_add comp1349(.out(wire1803), .cout(wire1804), .inA(wire1462), .inB(wire1464), .cin(wire1466));
	full_add comp1350(.out(wire1805), .cout(wire1806), .inA(wire1468), .inB(wire1470), .cin(wire1472));
	full_add comp1351(.out(wire1807), .cout(wire1808), .inA(wire1474), .inB(wire1475), .cin(wire1477));
	full_add comp1352(.out(wire1809), .cout(wire1810), .inA(wire1479), .inB(wire1481), .cin(wire1483));
	full_add comp1353(.out(wire1811), .cout(wire1812), .inA(wire913), .inB(wire944), .cin(wire975));
	full_add comp1354(.out(wire1813), .cout(wire1814), .inA(wire1006), .inB(wire1037), .cin(wire1068));
	full_add comp1355(.out(wire1815), .cout(wire1816), .inA(wire1099), .inB(wire1130), .cin(wire1476));
	full_add comp1356(.out(wire1817), .cout(wire1818), .inA(wire1478), .inB(wire1480), .cin(wire1482));
	full_add comp1357(.out(wire1819), .cout(wire1820), .inA(wire1484), .inB(wire1486), .cin(wire1487));
	full_add comp1358(.out(wire1821), .cout(wire1822), .inA(wire1489), .inB(wire1491), .cin(wire1493));
	full_add comp1359(.out(wire1823), .cout(wire1824), .inA(wire852), .inB(wire883), .cin(wire914));
	full_add comp1360(.out(wire1825), .cout(wire1826), .inA(wire945), .inB(wire976), .cin(wire1007));
	full_add comp1361(.out(wire1827), .cout(wire1828), .inA(wire1038), .inB(wire1069), .cin(wire1100));
	full_add comp1362(.out(wire1829), .cout(wire1830), .inA(wire1131), .inB(wire1488), .cin(wire1490));
	full_add comp1363(.out(wire1831), .cout(wire1832), .inA(wire1492), .inB(wire1494), .cin(wire1496));
	full_add comp1364(.out(wire1833), .cout(wire1834), .inA(wire1497), .inB(wire1499), .cin(wire1501));
	full_add comp1365(.out(wire1835), .cout(wire1836), .inA(wire791), .inB(wire822), .cin(wire853));
	full_add comp1366(.out(wire1837), .cout(wire1838), .inA(wire884), .inB(wire915), .cin(wire946));
	full_add comp1367(.out(wire1839), .cout(wire1840), .inA(wire977), .inB(wire1008), .cin(wire1039));
	full_add comp1368(.out(wire1841), .cout(wire1842), .inA(wire1070), .inB(wire1101), .cin(wire1132));
	full_add comp1369(.out(wire1843), .cout(wire1844), .inA(wire1498), .inB(wire1500), .cin(wire1502));
	full_add comp1370(.out(wire1845), .cout(wire1846), .inA(wire1504), .inB(wire1505), .cin(wire1507));
	full_add comp1371(.out(wire1847), .cout(wire1848), .inA(wire730), .inB(wire761), .cin(wire792));
	full_add comp1372(.out(wire1849), .cout(wire1850), .inA(wire823), .inB(wire854), .cin(wire885));
	full_add comp1373(.out(wire1851), .cout(wire1852), .inA(wire916), .inB(wire947), .cin(wire978));
	full_add comp1374(.out(wire1853), .cout(wire1854), .inA(wire1009), .inB(wire1040), .cin(wire1071));
	full_add comp1375(.out(wire1855), .cout(wire1856), .inA(wire1102), .inB(wire1133), .cin(wire1506));
	full_add comp1376(.out(wire1857), .cout(wire1858), .inA(wire1508), .inB(wire1510), .cin(wire1511));
	full_add comp1377(.out(wire1859), .cout(wire1860), .inA(wire669), .inB(wire700), .cin(wire731));
	full_add comp1378(.out(wire1861), .cout(wire1862), .inA(wire762), .inB(wire793), .cin(wire824));
	full_add comp1379(.out(wire1863), .cout(wire1864), .inA(wire855), .inB(wire886), .cin(wire917));
	full_add comp1380(.out(wire1865), .cout(wire1866), .inA(wire948), .inB(wire979), .cin(wire1010));
	full_add comp1381(.out(wire1867), .cout(wire1868), .inA(wire1041), .inB(wire1072), .cin(wire1103));
	full_add comp1382(.out(wire1869), .cout(wire1870), .inA(wire1134), .inB(wire1512), .cin(wire1514));
	full_add comp1383(.out(wire1871), .cout(wire1872), .inA(wire608), .inB(wire639), .cin(wire670));
	full_add comp1384(.out(wire1873), .cout(wire1874), .inA(wire701), .inB(wire732), .cin(wire763));
	full_add comp1385(.out(wire1875), .cout(wire1876), .inA(wire794), .inB(wire825), .cin(wire856));
	full_add comp1386(.out(wire1877), .cout(wire1878), .inA(wire887), .inB(wire918), .cin(wire949));
	full_add comp1387(.out(wire1879), .cout(wire1880), .inA(wire980), .inB(wire1011), .cin(wire1042));
	full_add comp1388(.out(wire1881), .cout(wire1882), .inA(wire1073), .inB(wire1104), .cin(wire1135));
	full_add comp1389(.out(wire1883), .cout(wire1884), .inA(wire640), .inB(wire671), .cin(wire702));
	full_add comp1390(.out(wire1885), .cout(wire1886), .inA(wire733), .inB(wire764), .cin(wire795));
	full_add comp1391(.out(wire1887), .cout(wire1888), .inA(wire826), .inB(wire857), .cin(wire888));
	full_add comp1392(.out(wire1889), .cout(wire1890), .inA(wire919), .inB(wire950), .cin(wire981));
	full_add comp1393(.out(wire1891), .cout(wire1892), .inA(wire1012), .inB(wire1043), .cin(wire1074));
	full_add comp1394(.out(wire1893), .cout(wire1894), .inA(wire672), .inB(wire703), .cin(wire734));
	full_add comp1395(.out(wire1895), .cout(wire1896), .inA(wire765), .inB(wire796), .cin(wire827));
	full_add comp1396(.out(wire1897), .cout(wire1898), .inA(wire858), .inB(wire889), .cin(wire920));
	full_add comp1397(.out(wire1899), .cout(wire1900), .inA(wire951), .inB(wire982), .cin(wire1013));
	full_add comp1398(.out(wire1901), .cout(wire1902), .inA(wire704), .inB(wire735), .cin(wire766));
	full_add comp1399(.out(wire1903), .cout(wire1904), .inA(wire797), .inB(wire828), .cin(wire859));
	full_add comp1400(.out(wire1905), .cout(wire1906), .inA(wire890), .inB(wire921), .cin(wire952));
	full_add comp1401(.out(wire1907), .cout(wire1908), .inA(wire736), .inB(wire767), .cin(wire798));
	full_add comp1402(.out(wire1909), .cout(wire1910), .inA(wire829), .inB(wire860), .cin(wire891));
	full_add comp1403(.out(wire1911), .cout(wire1912), .inA(wire768), .inB(wire799), .cin(wire830));
	half_add comp1404(.out(wire1913), .cout(wire1914), .inA(wire138), .inB(wire169));
	full_add comp1405(.out(wire1915), .cout(wire1916), .inA(wire139), .inB(wire170), .cin(wire201));
	half_add comp1406(.out(wire1917), .cout(wire1918), .inA(wire232), .inB(wire263));
	full_add comp1407(.out(wire1919), .cout(wire1920), .inA(wire140), .inB(wire171), .cin(wire202));
	full_add comp1408(.out(wire1921), .cout(wire1922), .inA(wire233), .inB(wire264), .cin(wire295));
	half_add comp1409(.out(wire1923), .cout(wire1924), .inA(wire326), .inB(wire357));
	full_add comp1410(.out(wire1925), .cout(wire1926), .inA(wire141), .inB(wire172), .cin(wire203));
	full_add comp1411(.out(wire1927), .cout(wire1928), .inA(wire234), .inB(wire265), .cin(wire296));
	full_add comp1412(.out(wire1929), .cout(wire1930), .inA(wire327), .inB(wire358), .cin(wire389));
	half_add comp1413(.out(wire1931), .cout(wire1932), .inA(wire420), .inB(wire451));
	full_add comp1414(.out(wire1933), .cout(wire1934), .inA(wire204), .inB(wire235), .cin(wire266));
	full_add comp1415(.out(wire1935), .cout(wire1936), .inA(wire297), .inB(wire328), .cin(wire359));
	full_add comp1416(.out(wire1937), .cout(wire1938), .inA(wire390), .inB(wire421), .cin(wire452));
	full_add comp1417(.out(wire1939), .cout(wire1940), .inA(wire483), .inB(wire514), .cin(wire545));
	full_add comp1418(.out(wire1941), .cout(wire1942), .inA(wire298), .inB(wire329), .cin(wire360));
	full_add comp1419(.out(wire1943), .cout(wire1944), .inA(wire391), .inB(wire422), .cin(wire453));
	full_add comp1420(.out(wire1945), .cout(wire1946), .inA(wire484), .inB(wire515), .cin(wire546));
	full_add comp1421(.out(wire1947), .cout(wire1948), .inA(wire577), .inB(wire1518), .cin(wire1519));
	full_add comp1422(.out(wire1949), .cout(wire1950), .inA(wire392), .inB(wire423), .cin(wire454));
	full_add comp1423(.out(wire1951), .cout(wire1952), .inA(wire485), .inB(wire516), .cin(wire547));
	full_add comp1424(.out(wire1953), .cout(wire1954), .inA(wire578), .inB(wire609), .cin(wire1520));
	full_add comp1425(.out(wire1955), .cout(wire1956), .inA(wire1522), .inB(wire1523), .cin(wire1525));
	full_add comp1426(.out(wire1957), .cout(wire1958), .inA(wire486), .inB(wire517), .cin(wire548));
	full_add comp1427(.out(wire1959), .cout(wire1960), .inA(wire579), .inB(wire610), .cin(wire641));
	full_add comp1428(.out(wire1961), .cout(wire1962), .inA(wire1524), .inB(wire1526), .cin(wire1528));
	full_add comp1429(.out(wire1963), .cout(wire1964), .inA(wire1529), .inB(wire1531), .cin(wire1533));
	full_add comp1430(.out(wire1965), .cout(wire1966), .inA(wire580), .inB(wire611), .cin(wire642));
	full_add comp1431(.out(wire1967), .cout(wire1968), .inA(wire673), .inB(wire1530), .cin(wire1532));
	full_add comp1432(.out(wire1969), .cout(wire1970), .inA(wire1534), .inB(wire1536), .cin(wire1537));
	full_add comp1433(.out(wire1971), .cout(wire1972), .inA(wire1539), .inB(wire1541), .cin(wire1543));
	full_add comp1434(.out(wire1973), .cout(wire1974), .inA(wire674), .inB(wire705), .cin(wire1538));
	full_add comp1435(.out(wire1975), .cout(wire1976), .inA(wire1540), .inB(wire1542), .cin(wire1544));
	full_add comp1436(.out(wire1977), .cout(wire1978), .inA(wire1546), .inB(wire1547), .cin(wire1549));
	full_add comp1437(.out(wire1979), .cout(wire1980), .inA(wire1551), .inB(wire1553), .cin(wire1555));
	full_add comp1438(.out(wire1981), .cout(wire1982), .inA(wire1193), .inB(wire1548), .cin(wire1550));
	full_add comp1439(.out(wire1983), .cout(wire1984), .inA(wire1552), .inB(wire1554), .cin(wire1556));
	full_add comp1440(.out(wire1985), .cout(wire1986), .inA(wire1558), .inB(wire1559), .cin(wire1561));
	full_add comp1441(.out(wire1987), .cout(wire1988), .inA(wire1563), .inB(wire1565), .cin(wire1567));
	full_add comp1442(.out(wire1989), .cout(wire1990), .inA(wire1197), .inB(wire1560), .cin(wire1562));
	full_add comp1443(.out(wire1991), .cout(wire1992), .inA(wire1564), .inB(wire1566), .cin(wire1568));
	full_add comp1444(.out(wire1993), .cout(wire1994), .inA(wire1570), .inB(wire1571), .cin(wire1573));
	full_add comp1445(.out(wire1995), .cout(wire1996), .inA(wire1575), .inB(wire1577), .cin(wire1579));
	full_add comp1446(.out(wire1997), .cout(wire1998), .inA(wire1203), .inB(wire1572), .cin(wire1574));
	full_add comp1447(.out(wire1999), .cout(wire2000), .inA(wire1576), .inB(wire1578), .cin(wire1580));
	full_add comp1448(.out(wire2001), .cout(wire2002), .inA(wire1582), .inB(wire1583), .cin(wire1585));
	full_add comp1449(.out(wire2003), .cout(wire2004), .inA(wire1587), .inB(wire1589), .cin(wire1591));
	full_add comp1450(.out(wire2005), .cout(wire2006), .inA(wire1211), .inB(wire1584), .cin(wire1586));
	full_add comp1451(.out(wire2007), .cout(wire2008), .inA(wire1588), .inB(wire1590), .cin(wire1592));
	full_add comp1452(.out(wire2009), .cout(wire2010), .inA(wire1594), .inB(wire1595), .cin(wire1597));
	full_add comp1453(.out(wire2011), .cout(wire2012), .inA(wire1599), .inB(wire1601), .cin(wire1603));
	full_add comp1454(.out(wire2013), .cout(wire2014), .inA(wire1221), .inB(wire1596), .cin(wire1598));
	full_add comp1455(.out(wire2015), .cout(wire2016), .inA(wire1600), .inB(wire1602), .cin(wire1604));
	full_add comp1456(.out(wire2017), .cout(wire2018), .inA(wire1606), .inB(wire1607), .cin(wire1609));
	full_add comp1457(.out(wire2019), .cout(wire2020), .inA(wire1611), .inB(wire1613), .cin(wire1615));
	full_add comp1458(.out(wire2021), .cout(wire2022), .inA(wire1233), .inB(wire1608), .cin(wire1610));
	full_add comp1459(.out(wire2023), .cout(wire2024), .inA(wire1612), .inB(wire1614), .cin(wire1616));
	full_add comp1460(.out(wire2025), .cout(wire2026), .inA(wire1618), .inB(wire1619), .cin(wire1621));
	full_add comp1461(.out(wire2027), .cout(wire2028), .inA(wire1623), .inB(wire1625), .cin(wire1627));
	full_add comp1462(.out(wire2029), .cout(wire2030), .inA(wire1247), .inB(wire1620), .cin(wire1622));
	full_add comp1463(.out(wire2031), .cout(wire2032), .inA(wire1624), .inB(wire1626), .cin(wire1628));
	full_add comp1464(.out(wire2033), .cout(wire2034), .inA(wire1630), .inB(wire1631), .cin(wire1633));
	full_add comp1465(.out(wire2035), .cout(wire2036), .inA(wire1635), .inB(wire1637), .cin(wire1639));
	full_add comp1466(.out(wire2037), .cout(wire2038), .inA(wire1263), .inB(wire1632), .cin(wire1634));
	full_add comp1467(.out(wire2039), .cout(wire2040), .inA(wire1636), .inB(wire1638), .cin(wire1640));
	full_add comp1468(.out(wire2041), .cout(wire2042), .inA(wire1642), .inB(wire1643), .cin(wire1645));
	full_add comp1469(.out(wire2043), .cout(wire2044), .inA(wire1647), .inB(wire1649), .cin(wire1651));
	full_add comp1470(.out(wire2045), .cout(wire2046), .inA(wire1281), .inB(wire1644), .cin(wire1646));
	full_add comp1471(.out(wire2047), .cout(wire2048), .inA(wire1648), .inB(wire1650), .cin(wire1652));
	full_add comp1472(.out(wire2049), .cout(wire2050), .inA(wire1654), .inB(wire1655), .cin(wire1657));
	full_add comp1473(.out(wire2051), .cout(wire2052), .inA(wire1659), .inB(wire1661), .cin(wire1663));
	full_add comp1474(.out(wire2053), .cout(wire2054), .inA(wire1299), .inB(wire1656), .cin(wire1658));
	full_add comp1475(.out(wire2055), .cout(wire2056), .inA(wire1660), .inB(wire1662), .cin(wire1664));
	full_add comp1476(.out(wire2057), .cout(wire2058), .inA(wire1666), .inB(wire1667), .cin(wire1669));
	full_add comp1477(.out(wire2059), .cout(wire2060), .inA(wire1671), .inB(wire1673), .cin(wire1675));
	full_add comp1478(.out(wire2061), .cout(wire2062), .inA(wire1317), .inB(wire1668), .cin(wire1670));
	full_add comp1479(.out(wire2063), .cout(wire2064), .inA(wire1672), .inB(wire1674), .cin(wire1676));
	full_add comp1480(.out(wire2065), .cout(wire2066), .inA(wire1678), .inB(wire1679), .cin(wire1681));
	full_add comp1481(.out(wire2067), .cout(wire2068), .inA(wire1683), .inB(wire1685), .cin(wire1687));
	full_add comp1482(.out(wire2069), .cout(wire2070), .inA(wire1335), .inB(wire1680), .cin(wire1682));
	full_add comp1483(.out(wire2071), .cout(wire2072), .inA(wire1684), .inB(wire1686), .cin(wire1688));
	full_add comp1484(.out(wire2073), .cout(wire2074), .inA(wire1690), .inB(wire1691), .cin(wire1693));
	full_add comp1485(.out(wire2075), .cout(wire2076), .inA(wire1695), .inB(wire1697), .cin(wire1699));
	full_add comp1486(.out(wire2077), .cout(wire2078), .inA(wire1353), .inB(wire1692), .cin(wire1694));
	full_add comp1487(.out(wire2079), .cout(wire2080), .inA(wire1696), .inB(wire1698), .cin(wire1700));
	full_add comp1488(.out(wire2081), .cout(wire2082), .inA(wire1702), .inB(wire1703), .cin(wire1705));
	full_add comp1489(.out(wire2083), .cout(wire2084), .inA(wire1707), .inB(wire1709), .cin(wire1711));
	full_add comp1490(.out(wire2085), .cout(wire2086), .inA(wire1371), .inB(wire1704), .cin(wire1706));
	full_add comp1491(.out(wire2087), .cout(wire2088), .inA(wire1708), .inB(wire1710), .cin(wire1712));
	full_add comp1492(.out(wire2089), .cout(wire2090), .inA(wire1714), .inB(wire1715), .cin(wire1717));
	full_add comp1493(.out(wire2091), .cout(wire2092), .inA(wire1719), .inB(wire1721), .cin(wire1723));
	full_add comp1494(.out(wire2093), .cout(wire2094), .inA(wire1389), .inB(wire1716), .cin(wire1718));
	full_add comp1495(.out(wire2095), .cout(wire2096), .inA(wire1720), .inB(wire1722), .cin(wire1724));
	full_add comp1496(.out(wire2097), .cout(wire2098), .inA(wire1726), .inB(wire1727), .cin(wire1729));
	full_add comp1497(.out(wire2099), .cout(wire2100), .inA(wire1731), .inB(wire1733), .cin(wire1735));
	full_add comp1498(.out(wire2101), .cout(wire2102), .inA(wire1407), .inB(wire1728), .cin(wire1730));
	full_add comp1499(.out(wire2103), .cout(wire2104), .inA(wire1732), .inB(wire1734), .cin(wire1736));
	full_add comp1500(.out(wire2105), .cout(wire2106), .inA(wire1738), .inB(wire1739), .cin(wire1741));
	full_add comp1501(.out(wire2107), .cout(wire2108), .inA(wire1743), .inB(wire1745), .cin(wire1747));
	full_add comp1502(.out(wire2109), .cout(wire2110), .inA(wire1425), .inB(wire1740), .cin(wire1742));
	full_add comp1503(.out(wire2111), .cout(wire2112), .inA(wire1744), .inB(wire1746), .cin(wire1748));
	full_add comp1504(.out(wire2113), .cout(wire2114), .inA(wire1750), .inB(wire1751), .cin(wire1753));
	full_add comp1505(.out(wire2115), .cout(wire2116), .inA(wire1755), .inB(wire1757), .cin(wire1759));
	full_add comp1506(.out(wire2117), .cout(wire2118), .inA(wire1443), .inB(wire1752), .cin(wire1754));
	full_add comp1507(.out(wire2119), .cout(wire2120), .inA(wire1756), .inB(wire1758), .cin(wire1760));
	full_add comp1508(.out(wire2121), .cout(wire2122), .inA(wire1762), .inB(wire1763), .cin(wire1765));
	full_add comp1509(.out(wire2123), .cout(wire2124), .inA(wire1767), .inB(wire1769), .cin(wire1771));
	full_add comp1510(.out(wire2125), .cout(wire2126), .inA(wire1459), .inB(wire1764), .cin(wire1766));
	full_add comp1511(.out(wire2127), .cout(wire2128), .inA(wire1768), .inB(wire1770), .cin(wire1772));
	full_add comp1512(.out(wire2129), .cout(wire2130), .inA(wire1774), .inB(wire1775), .cin(wire1777));
	full_add comp1513(.out(wire2131), .cout(wire2132), .inA(wire1779), .inB(wire1781), .cin(wire1783));
	full_add comp1514(.out(wire2133), .cout(wire2134), .inA(wire1473), .inB(wire1776), .cin(wire1778));
	full_add comp1515(.out(wire2135), .cout(wire2136), .inA(wire1780), .inB(wire1782), .cin(wire1784));
	full_add comp1516(.out(wire2137), .cout(wire2138), .inA(wire1786), .inB(wire1787), .cin(wire1789));
	full_add comp1517(.out(wire2139), .cout(wire2140), .inA(wire1791), .inB(wire1793), .cin(wire1795));
	full_add comp1518(.out(wire2141), .cout(wire2142), .inA(wire1485), .inB(wire1788), .cin(wire1790));
	full_add comp1519(.out(wire2143), .cout(wire2144), .inA(wire1792), .inB(wire1794), .cin(wire1796));
	full_add comp1520(.out(wire2145), .cout(wire2146), .inA(wire1798), .inB(wire1799), .cin(wire1801));
	full_add comp1521(.out(wire2147), .cout(wire2148), .inA(wire1803), .inB(wire1805), .cin(wire1807));
	full_add comp1522(.out(wire2149), .cout(wire2150), .inA(wire1495), .inB(wire1800), .cin(wire1802));
	full_add comp1523(.out(wire2151), .cout(wire2152), .inA(wire1804), .inB(wire1806), .cin(wire1808));
	full_add comp1524(.out(wire2153), .cout(wire2154), .inA(wire1810), .inB(wire1811), .cin(wire1813));
	full_add comp1525(.out(wire2155), .cout(wire2156), .inA(wire1815), .inB(wire1817), .cin(wire1819));
	full_add comp1526(.out(wire2157), .cout(wire2158), .inA(wire1503), .inB(wire1812), .cin(wire1814));
	full_add comp1527(.out(wire2159), .cout(wire2160), .inA(wire1816), .inB(wire1818), .cin(wire1820));
	full_add comp1528(.out(wire2161), .cout(wire2162), .inA(wire1822), .inB(wire1823), .cin(wire1825));
	full_add comp1529(.out(wire2163), .cout(wire2164), .inA(wire1827), .inB(wire1829), .cin(wire1831));
	full_add comp1530(.out(wire2165), .cout(wire2166), .inA(wire1509), .inB(wire1824), .cin(wire1826));
	full_add comp1531(.out(wire2167), .cout(wire2168), .inA(wire1828), .inB(wire1830), .cin(wire1832));
	full_add comp1532(.out(wire2169), .cout(wire2170), .inA(wire1834), .inB(wire1835), .cin(wire1837));
	full_add comp1533(.out(wire2171), .cout(wire2172), .inA(wire1839), .inB(wire1841), .cin(wire1843));
	full_add comp1534(.out(wire2173), .cout(wire2174), .inA(wire1513), .inB(wire1836), .cin(wire1838));
	full_add comp1535(.out(wire2175), .cout(wire2176), .inA(wire1840), .inB(wire1842), .cin(wire1844));
	full_add comp1536(.out(wire2177), .cout(wire2178), .inA(wire1846), .inB(wire1847), .cin(wire1849));
	full_add comp1537(.out(wire2179), .cout(wire2180), .inA(wire1851), .inB(wire1853), .cin(wire1855));
	full_add comp1538(.out(wire2181), .cout(wire2182), .inA(wire1515), .inB(wire1848), .cin(wire1850));
	full_add comp1539(.out(wire2183), .cout(wire2184), .inA(wire1852), .inB(wire1854), .cin(wire1856));
	full_add comp1540(.out(wire2185), .cout(wire2186), .inA(wire1858), .inB(wire1859), .cin(wire1861));
	full_add comp1541(.out(wire2187), .cout(wire2188), .inA(wire1863), .inB(wire1865), .cin(wire1867));
	full_add comp1542(.out(wire2189), .cout(wire2190), .inA(wire1516), .inB(wire1860), .cin(wire1862));
	full_add comp1543(.out(wire2191), .cout(wire2192), .inA(wire1864), .inB(wire1866), .cin(wire1868));
	full_add comp1544(.out(wire2193), .cout(wire2194), .inA(wire1870), .inB(wire1871), .cin(wire1873));
	full_add comp1545(.out(wire2195), .cout(wire2196), .inA(wire1875), .inB(wire1877), .cin(wire1879));
	full_add comp1546(.out(wire2197), .cout(wire2198), .inA(wire1105), .inB(wire1136), .cin(wire1872));
	full_add comp1547(.out(wire2199), .cout(wire2200), .inA(wire1874), .inB(wire1876), .cin(wire1878));
	full_add comp1548(.out(wire2201), .cout(wire2202), .inA(wire1880), .inB(wire1882), .cin(wire1883));
	full_add comp1549(.out(wire2203), .cout(wire2204), .inA(wire1885), .inB(wire1887), .cin(wire1889));
	full_add comp1550(.out(wire2205), .cout(wire2206), .inA(wire1044), .inB(wire1075), .cin(wire1106));
	full_add comp1551(.out(wire2207), .cout(wire2208), .inA(wire1137), .inB(wire1884), .cin(wire1886));
	full_add comp1552(.out(wire2209), .cout(wire2210), .inA(wire1888), .inB(wire1890), .cin(wire1892));
	full_add comp1553(.out(wire2211), .cout(wire2212), .inA(wire1893), .inB(wire1895), .cin(wire1897));
	full_add comp1554(.out(wire2213), .cout(wire2214), .inA(wire983), .inB(wire1014), .cin(wire1045));
	full_add comp1555(.out(wire2215), .cout(wire2216), .inA(wire1076), .inB(wire1107), .cin(wire1138));
	full_add comp1556(.out(wire2217), .cout(wire2218), .inA(wire1894), .inB(wire1896), .cin(wire1898));
	full_add comp1557(.out(wire2219), .cout(wire2220), .inA(wire1900), .inB(wire1901), .cin(wire1903));
	full_add comp1558(.out(wire2221), .cout(wire2222), .inA(wire922), .inB(wire953), .cin(wire984));
	full_add comp1559(.out(wire2223), .cout(wire2224), .inA(wire1015), .inB(wire1046), .cin(wire1077));
	full_add comp1560(.out(wire2225), .cout(wire2226), .inA(wire1108), .inB(wire1139), .cin(wire1902));
	full_add comp1561(.out(wire2227), .cout(wire2228), .inA(wire1904), .inB(wire1906), .cin(wire1907));
	full_add comp1562(.out(wire2229), .cout(wire2230), .inA(wire861), .inB(wire892), .cin(wire923));
	full_add comp1563(.out(wire2231), .cout(wire2232), .inA(wire954), .inB(wire985), .cin(wire1016));
	full_add comp1564(.out(wire2233), .cout(wire2234), .inA(wire1047), .inB(wire1078), .cin(wire1109));
	full_add comp1565(.out(wire2235), .cout(wire2236), .inA(wire1140), .inB(wire1908), .cin(wire1910));
	full_add comp1566(.out(wire2237), .cout(wire2238), .inA(wire800), .inB(wire831), .cin(wire862));
	full_add comp1567(.out(wire2239), .cout(wire2240), .inA(wire893), .inB(wire924), .cin(wire955));
	full_add comp1568(.out(wire2241), .cout(wire2242), .inA(wire986), .inB(wire1017), .cin(wire1048));
	full_add comp1569(.out(wire2243), .cout(wire2244), .inA(wire1079), .inB(wire1110), .cin(wire1141));
	full_add comp1570(.out(wire2245), .cout(wire2246), .inA(wire832), .inB(wire863), .cin(wire894));
	full_add comp1571(.out(wire2247), .cout(wire2248), .inA(wire925), .inB(wire956), .cin(wire987));
	full_add comp1572(.out(wire2249), .cout(wire2250), .inA(wire1018), .inB(wire1049), .cin(wire1080));
	full_add comp1573(.out(wire2251), .cout(wire2252), .inA(wire864), .inB(wire895), .cin(wire926));
	full_add comp1574(.out(wire2253), .cout(wire2254), .inA(wire957), .inB(wire988), .cin(wire1019));
	full_add comp1575(.out(wire2255), .cout(wire2256), .inA(wire896), .inB(wire927), .cin(wire958));
	half_add comp1576(.out(wire2257), .cout(wire2258), .inA(wire135), .inB(wire166));
	full_add comp1577(.out(wire2259), .cout(wire2260), .inA(wire136), .inB(wire167), .cin(wire198));
	half_add comp1578(.out(wire2261), .cout(wire2262), .inA(wire229), .inB(wire260));
	full_add comp1579(.out(wire2263), .cout(wire2264), .inA(wire137), .inB(wire168), .cin(wire199));
	full_add comp1580(.out(wire2265), .cout(wire2266), .inA(wire230), .inB(wire261), .cin(wire292));
	half_add comp1581(.out(wire2267), .cout(wire2268), .inA(wire323), .inB(wire354));
	full_add comp1582(.out(wire2269), .cout(wire2270), .inA(wire200), .inB(wire231), .cin(wire262));
	full_add comp1583(.out(wire2271), .cout(wire2272), .inA(wire293), .inB(wire324), .cin(wire355));
	full_add comp1584(.out(wire2273), .cout(wire2274), .inA(wire386), .inB(wire417), .cin(wire1913));
	full_add comp1585(.out(wire2275), .cout(wire2276), .inA(wire294), .inB(wire325), .cin(wire356));
	full_add comp1586(.out(wire2277), .cout(wire2278), .inA(wire387), .inB(wire418), .cin(wire449));
	full_add comp1587(.out(wire2279), .cout(wire2280), .inA(wire1914), .inB(wire1915), .cin(wire1917));
	full_add comp1588(.out(wire2281), .cout(wire2282), .inA(wire388), .inB(wire419), .cin(wire450));
	full_add comp1589(.out(wire2283), .cout(wire2284), .inA(wire481), .inB(wire1916), .cin(wire1918));
	full_add comp1590(.out(wire2285), .cout(wire2286), .inA(wire1919), .inB(wire1921), .cin(wire1923));
	full_add comp1591(.out(wire2287), .cout(wire2288), .inA(wire482), .inB(wire513), .cin(wire1920));
	full_add comp1592(.out(wire2289), .cout(wire2290), .inA(wire1922), .inB(wire1924), .cin(wire1925));
	full_add comp1593(.out(wire2291), .cout(wire2292), .inA(wire1927), .inB(wire1929), .cin(wire1931));
	full_add comp1594(.out(wire2293), .cout(wire2294), .inA(wire1517), .inB(wire1926), .cin(wire1928));
	full_add comp1595(.out(wire2295), .cout(wire2296), .inA(wire1930), .inB(wire1932), .cin(wire1933));
	full_add comp1596(.out(wire2297), .cout(wire2298), .inA(wire1935), .inB(wire1937), .cin(wire1939));
	full_add comp1597(.out(wire2299), .cout(wire2300), .inA(wire1521), .inB(wire1934), .cin(wire1936));
	full_add comp1598(.out(wire2301), .cout(wire2302), .inA(wire1938), .inB(wire1940), .cin(wire1941));
	full_add comp1599(.out(wire2303), .cout(wire2304), .inA(wire1943), .inB(wire1945), .cin(wire1947));
	full_add comp1600(.out(wire2305), .cout(wire2306), .inA(wire1527), .inB(wire1942), .cin(wire1944));
	full_add comp1601(.out(wire2307), .cout(wire2308), .inA(wire1946), .inB(wire1948), .cin(wire1949));
	full_add comp1602(.out(wire2309), .cout(wire2310), .inA(wire1951), .inB(wire1953), .cin(wire1955));
	full_add comp1603(.out(wire2311), .cout(wire2312), .inA(wire1535), .inB(wire1950), .cin(wire1952));
	full_add comp1604(.out(wire2313), .cout(wire2314), .inA(wire1954), .inB(wire1956), .cin(wire1957));
	full_add comp1605(.out(wire2315), .cout(wire2316), .inA(wire1959), .inB(wire1961), .cin(wire1963));
	full_add comp1606(.out(wire2317), .cout(wire2318), .inA(wire1545), .inB(wire1958), .cin(wire1960));
	full_add comp1607(.out(wire2319), .cout(wire2320), .inA(wire1962), .inB(wire1964), .cin(wire1965));
	full_add comp1608(.out(wire2321), .cout(wire2322), .inA(wire1967), .inB(wire1969), .cin(wire1971));
	full_add comp1609(.out(wire2323), .cout(wire2324), .inA(wire1557), .inB(wire1966), .cin(wire1968));
	full_add comp1610(.out(wire2325), .cout(wire2326), .inA(wire1970), .inB(wire1972), .cin(wire1973));
	full_add comp1611(.out(wire2327), .cout(wire2328), .inA(wire1975), .inB(wire1977), .cin(wire1979));
	full_add comp1612(.out(wire2329), .cout(wire2330), .inA(wire1569), .inB(wire1974), .cin(wire1976));
	full_add comp1613(.out(wire2331), .cout(wire2332), .inA(wire1978), .inB(wire1980), .cin(wire1981));
	full_add comp1614(.out(wire2333), .cout(wire2334), .inA(wire1983), .inB(wire1985), .cin(wire1987));
	full_add comp1615(.out(wire2335), .cout(wire2336), .inA(wire1581), .inB(wire1982), .cin(wire1984));
	full_add comp1616(.out(wire2337), .cout(wire2338), .inA(wire1986), .inB(wire1988), .cin(wire1989));
	full_add comp1617(.out(wire2339), .cout(wire2340), .inA(wire1991), .inB(wire1993), .cin(wire1995));
	full_add comp1618(.out(wire2341), .cout(wire2342), .inA(wire1593), .inB(wire1990), .cin(wire1992));
	full_add comp1619(.out(wire2343), .cout(wire2344), .inA(wire1994), .inB(wire1996), .cin(wire1997));
	full_add comp1620(.out(wire2345), .cout(wire2346), .inA(wire1999), .inB(wire2001), .cin(wire2003));
	full_add comp1621(.out(wire2347), .cout(wire2348), .inA(wire1605), .inB(wire1998), .cin(wire2000));
	full_add comp1622(.out(wire2349), .cout(wire2350), .inA(wire2002), .inB(wire2004), .cin(wire2005));
	full_add comp1623(.out(wire2351), .cout(wire2352), .inA(wire2007), .inB(wire2009), .cin(wire2011));
	full_add comp1624(.out(wire2353), .cout(wire2354), .inA(wire1617), .inB(wire2006), .cin(wire2008));
	full_add comp1625(.out(wire2355), .cout(wire2356), .inA(wire2010), .inB(wire2012), .cin(wire2013));
	full_add comp1626(.out(wire2357), .cout(wire2358), .inA(wire2015), .inB(wire2017), .cin(wire2019));
	full_add comp1627(.out(wire2359), .cout(wire2360), .inA(wire1629), .inB(wire2014), .cin(wire2016));
	full_add comp1628(.out(wire2361), .cout(wire2362), .inA(wire2018), .inB(wire2020), .cin(wire2021));
	full_add comp1629(.out(wire2363), .cout(wire2364), .inA(wire2023), .inB(wire2025), .cin(wire2027));
	full_add comp1630(.out(wire2365), .cout(wire2366), .inA(wire1641), .inB(wire2022), .cin(wire2024));
	full_add comp1631(.out(wire2367), .cout(wire2368), .inA(wire2026), .inB(wire2028), .cin(wire2029));
	full_add comp1632(.out(wire2369), .cout(wire2370), .inA(wire2031), .inB(wire2033), .cin(wire2035));
	full_add comp1633(.out(wire2371), .cout(wire2372), .inA(wire1653), .inB(wire2030), .cin(wire2032));
	full_add comp1634(.out(wire2373), .cout(wire2374), .inA(wire2034), .inB(wire2036), .cin(wire2037));
	full_add comp1635(.out(wire2375), .cout(wire2376), .inA(wire2039), .inB(wire2041), .cin(wire2043));
	full_add comp1636(.out(wire2377), .cout(wire2378), .inA(wire1665), .inB(wire2038), .cin(wire2040));
	full_add comp1637(.out(wire2379), .cout(wire2380), .inA(wire2042), .inB(wire2044), .cin(wire2045));
	full_add comp1638(.out(wire2381), .cout(wire2382), .inA(wire2047), .inB(wire2049), .cin(wire2051));
	full_add comp1639(.out(wire2383), .cout(wire2384), .inA(wire1677), .inB(wire2046), .cin(wire2048));
	full_add comp1640(.out(wire2385), .cout(wire2386), .inA(wire2050), .inB(wire2052), .cin(wire2053));
	full_add comp1641(.out(wire2387), .cout(wire2388), .inA(wire2055), .inB(wire2057), .cin(wire2059));
	full_add comp1642(.out(wire2389), .cout(wire2390), .inA(wire1689), .inB(wire2054), .cin(wire2056));
	full_add comp1643(.out(wire2391), .cout(wire2392), .inA(wire2058), .inB(wire2060), .cin(wire2061));
	full_add comp1644(.out(wire2393), .cout(wire2394), .inA(wire2063), .inB(wire2065), .cin(wire2067));
	full_add comp1645(.out(wire2395), .cout(wire2396), .inA(wire1701), .inB(wire2062), .cin(wire2064));
	full_add comp1646(.out(wire2397), .cout(wire2398), .inA(wire2066), .inB(wire2068), .cin(wire2069));
	full_add comp1647(.out(wire2399), .cout(wire2400), .inA(wire2071), .inB(wire2073), .cin(wire2075));
	full_add comp1648(.out(wire2401), .cout(wire2402), .inA(wire1713), .inB(wire2070), .cin(wire2072));
	full_add comp1649(.out(wire2403), .cout(wire2404), .inA(wire2074), .inB(wire2076), .cin(wire2077));
	full_add comp1650(.out(wire2405), .cout(wire2406), .inA(wire2079), .inB(wire2081), .cin(wire2083));
	full_add comp1651(.out(wire2407), .cout(wire2408), .inA(wire1725), .inB(wire2078), .cin(wire2080));
	full_add comp1652(.out(wire2409), .cout(wire2410), .inA(wire2082), .inB(wire2084), .cin(wire2085));
	full_add comp1653(.out(wire2411), .cout(wire2412), .inA(wire2087), .inB(wire2089), .cin(wire2091));
	full_add comp1654(.out(wire2413), .cout(wire2414), .inA(wire1737), .inB(wire2086), .cin(wire2088));
	full_add comp1655(.out(wire2415), .cout(wire2416), .inA(wire2090), .inB(wire2092), .cin(wire2093));
	full_add comp1656(.out(wire2417), .cout(wire2418), .inA(wire2095), .inB(wire2097), .cin(wire2099));
	full_add comp1657(.out(wire2419), .cout(wire2420), .inA(wire1749), .inB(wire2094), .cin(wire2096));
	full_add comp1658(.out(wire2421), .cout(wire2422), .inA(wire2098), .inB(wire2100), .cin(wire2101));
	full_add comp1659(.out(wire2423), .cout(wire2424), .inA(wire2103), .inB(wire2105), .cin(wire2107));
	full_add comp1660(.out(wire2425), .cout(wire2426), .inA(wire1761), .inB(wire2102), .cin(wire2104));
	full_add comp1661(.out(wire2427), .cout(wire2428), .inA(wire2106), .inB(wire2108), .cin(wire2109));
	full_add comp1662(.out(wire2429), .cout(wire2430), .inA(wire2111), .inB(wire2113), .cin(wire2115));
	full_add comp1663(.out(wire2431), .cout(wire2432), .inA(wire1773), .inB(wire2110), .cin(wire2112));
	full_add comp1664(.out(wire2433), .cout(wire2434), .inA(wire2114), .inB(wire2116), .cin(wire2117));
	full_add comp1665(.out(wire2435), .cout(wire2436), .inA(wire2119), .inB(wire2121), .cin(wire2123));
	full_add comp1666(.out(wire2437), .cout(wire2438), .inA(wire1785), .inB(wire2118), .cin(wire2120));
	full_add comp1667(.out(wire2439), .cout(wire2440), .inA(wire2122), .inB(wire2124), .cin(wire2125));
	full_add comp1668(.out(wire2441), .cout(wire2442), .inA(wire2127), .inB(wire2129), .cin(wire2131));
	full_add comp1669(.out(wire2443), .cout(wire2444), .inA(wire1797), .inB(wire2126), .cin(wire2128));
	full_add comp1670(.out(wire2445), .cout(wire2446), .inA(wire2130), .inB(wire2132), .cin(wire2133));
	full_add comp1671(.out(wire2447), .cout(wire2448), .inA(wire2135), .inB(wire2137), .cin(wire2139));
	full_add comp1672(.out(wire2449), .cout(wire2450), .inA(wire1809), .inB(wire2134), .cin(wire2136));
	full_add comp1673(.out(wire2451), .cout(wire2452), .inA(wire2138), .inB(wire2140), .cin(wire2141));
	full_add comp1674(.out(wire2453), .cout(wire2454), .inA(wire2143), .inB(wire2145), .cin(wire2147));
	full_add comp1675(.out(wire2455), .cout(wire2456), .inA(wire1821), .inB(wire2142), .cin(wire2144));
	full_add comp1676(.out(wire2457), .cout(wire2458), .inA(wire2146), .inB(wire2148), .cin(wire2149));
	full_add comp1677(.out(wire2459), .cout(wire2460), .inA(wire2151), .inB(wire2153), .cin(wire2155));
	full_add comp1678(.out(wire2461), .cout(wire2462), .inA(wire1833), .inB(wire2150), .cin(wire2152));
	full_add comp1679(.out(wire2463), .cout(wire2464), .inA(wire2154), .inB(wire2156), .cin(wire2157));
	full_add comp1680(.out(wire2465), .cout(wire2466), .inA(wire2159), .inB(wire2161), .cin(wire2163));
	full_add comp1681(.out(wire2467), .cout(wire2468), .inA(wire1845), .inB(wire2158), .cin(wire2160));
	full_add comp1682(.out(wire2469), .cout(wire2470), .inA(wire2162), .inB(wire2164), .cin(wire2165));
	full_add comp1683(.out(wire2471), .cout(wire2472), .inA(wire2167), .inB(wire2169), .cin(wire2171));
	full_add comp1684(.out(wire2473), .cout(wire2474), .inA(wire1857), .inB(wire2166), .cin(wire2168));
	full_add comp1685(.out(wire2475), .cout(wire2476), .inA(wire2170), .inB(wire2172), .cin(wire2173));
	full_add comp1686(.out(wire2477), .cout(wire2478), .inA(wire2175), .inB(wire2177), .cin(wire2179));
	full_add comp1687(.out(wire2479), .cout(wire2480), .inA(wire1869), .inB(wire2174), .cin(wire2176));
	full_add comp1688(.out(wire2481), .cout(wire2482), .inA(wire2178), .inB(wire2180), .cin(wire2181));
	full_add comp1689(.out(wire2483), .cout(wire2484), .inA(wire2183), .inB(wire2185), .cin(wire2187));
	full_add comp1690(.out(wire2485), .cout(wire2486), .inA(wire1881), .inB(wire2182), .cin(wire2184));
	full_add comp1691(.out(wire2487), .cout(wire2488), .inA(wire2186), .inB(wire2188), .cin(wire2189));
	full_add comp1692(.out(wire2489), .cout(wire2490), .inA(wire2191), .inB(wire2193), .cin(wire2195));
	full_add comp1693(.out(wire2491), .cout(wire2492), .inA(wire1891), .inB(wire2190), .cin(wire2192));
	full_add comp1694(.out(wire2493), .cout(wire2494), .inA(wire2194), .inB(wire2196), .cin(wire2197));
	full_add comp1695(.out(wire2495), .cout(wire2496), .inA(wire2199), .inB(wire2201), .cin(wire2203));
	full_add comp1696(.out(wire2497), .cout(wire2498), .inA(wire1899), .inB(wire2198), .cin(wire2200));
	full_add comp1697(.out(wire2499), .cout(wire2500), .inA(wire2202), .inB(wire2204), .cin(wire2205));
	full_add comp1698(.out(wire2501), .cout(wire2502), .inA(wire2207), .inB(wire2209), .cin(wire2211));
	full_add comp1699(.out(wire2503), .cout(wire2504), .inA(wire1905), .inB(wire2206), .cin(wire2208));
	full_add comp1700(.out(wire2505), .cout(wire2506), .inA(wire2210), .inB(wire2212), .cin(wire2213));
	full_add comp1701(.out(wire2507), .cout(wire2508), .inA(wire2215), .inB(wire2217), .cin(wire2219));
	full_add comp1702(.out(wire2509), .cout(wire2510), .inA(wire1909), .inB(wire2214), .cin(wire2216));
	full_add comp1703(.out(wire2511), .cout(wire2512), .inA(wire2218), .inB(wire2220), .cin(wire2221));
	full_add comp1704(.out(wire2513), .cout(wire2514), .inA(wire2223), .inB(wire2225), .cin(wire2227));
	full_add comp1705(.out(wire2515), .cout(wire2516), .inA(wire1911), .inB(wire2222), .cin(wire2224));
	full_add comp1706(.out(wire2517), .cout(wire2518), .inA(wire2226), .inB(wire2228), .cin(wire2229));
	full_add comp1707(.out(wire2519), .cout(wire2520), .inA(wire2231), .inB(wire2233), .cin(wire2235));
	full_add comp1708(.out(wire2521), .cout(wire2522), .inA(wire1912), .inB(wire2230), .cin(wire2232));
	full_add comp1709(.out(wire2523), .cout(wire2524), .inA(wire2234), .inB(wire2236), .cin(wire2237));
	full_add comp1710(.out(wire2525), .cout(wire2526), .inA(wire2239), .inB(wire2241), .cin(wire2243));
	full_add comp1711(.out(wire2527), .cout(wire2528), .inA(wire1111), .inB(wire1142), .cin(wire2238));
	full_add comp1712(.out(wire2529), .cout(wire2530), .inA(wire2240), .inB(wire2242), .cin(wire2244));
	full_add comp1713(.out(wire2531), .cout(wire2532), .inA(wire2245), .inB(wire2247), .cin(wire2249));
	full_add comp1714(.out(wire2533), .cout(wire2534), .inA(wire1050), .inB(wire1081), .cin(wire1112));
	full_add comp1715(.out(wire2535), .cout(wire2536), .inA(wire1143), .inB(wire2246), .cin(wire2248));
	full_add comp1716(.out(wire2537), .cout(wire2538), .inA(wire2250), .inB(wire2251), .cin(wire2253));
	full_add comp1717(.out(wire2539), .cout(wire2540), .inA(wire989), .inB(wire1020), .cin(wire1051));
	full_add comp1718(.out(wire2541), .cout(wire2542), .inA(wire1082), .inB(wire1113), .cin(wire1144));
	full_add comp1719(.out(wire2543), .cout(wire2544), .inA(wire2252), .inB(wire2254), .cin(wire2255));
	full_add comp1720(.out(wire2545), .cout(wire2546), .inA(wire928), .inB(wire959), .cin(wire990));
	full_add comp1721(.out(wire2547), .cout(wire2548), .inA(wire1021), .inB(wire1052), .cin(wire1083));
	full_add comp1722(.out(wire2549), .cout(wire2550), .inA(wire1114), .inB(wire1145), .cin(wire2256));
	full_add comp1723(.out(wire2551), .cout(wire2552), .inA(wire960), .inB(wire991), .cin(wire1022));
	full_add comp1724(.out(wire2553), .cout(wire2554), .inA(wire1053), .inB(wire1084), .cin(wire1115));
	full_add comp1725(.out(wire2555), .cout(wire2556), .inA(wire992), .inB(wire1023), .cin(wire1054));
	half_add comp1726(.out(wire2557), .cout(wire2558), .inA(wire133), .inB(wire164));
	full_add comp1727(.out(wire2559), .cout(wire2560), .inA(wire134), .inB(wire165), .cin(wire196));
	half_add comp1728(.out(wire2561), .cout(wire2562), .inA(wire227), .inB(wire258));
	full_add comp1729(.out(wire2563), .cout(wire2564), .inA(wire197), .inB(wire228), .cin(wire259));
	full_add comp1730(.out(wire2565), .cout(wire2566), .inA(wire290), .inB(wire321), .cin(wire2257));
	full_add comp1731(.out(wire2567), .cout(wire2568), .inA(wire291), .inB(wire322), .cin(wire353));
	full_add comp1732(.out(wire2569), .cout(wire2570), .inA(wire2258), .inB(wire2259), .cin(wire2261));
	full_add comp1733(.out(wire2571), .cout(wire2572), .inA(wire385), .inB(wire2260), .cin(wire2262));
	full_add comp1734(.out(wire2573), .cout(wire2574), .inA(wire2263), .inB(wire2265), .cin(wire2267));
	full_add comp1735(.out(wire2575), .cout(wire2576), .inA(wire2264), .inB(wire2266), .cin(wire2268));
	full_add comp1736(.out(wire2577), .cout(wire2578), .inA(wire2269), .inB(wire2271), .cin(wire2273));
	full_add comp1737(.out(wire2579), .cout(wire2580), .inA(wire2270), .inB(wire2272), .cin(wire2274));
	full_add comp1738(.out(wire2581), .cout(wire2582), .inA(wire2275), .inB(wire2277), .cin(wire2279));
	full_add comp1739(.out(wire2583), .cout(wire2584), .inA(wire2276), .inB(wire2278), .cin(wire2280));
	full_add comp1740(.out(wire2585), .cout(wire2586), .inA(wire2281), .inB(wire2283), .cin(wire2285));
	full_add comp1741(.out(wire2587), .cout(wire2588), .inA(wire2282), .inB(wire2284), .cin(wire2286));
	full_add comp1742(.out(wire2589), .cout(wire2590), .inA(wire2287), .inB(wire2289), .cin(wire2291));
	full_add comp1743(.out(wire2591), .cout(wire2592), .inA(wire2288), .inB(wire2290), .cin(wire2292));
	full_add comp1744(.out(wire2593), .cout(wire2594), .inA(wire2293), .inB(wire2295), .cin(wire2297));
	full_add comp1745(.out(wire2595), .cout(wire2596), .inA(wire2294), .inB(wire2296), .cin(wire2298));
	full_add comp1746(.out(wire2597), .cout(wire2598), .inA(wire2299), .inB(wire2301), .cin(wire2303));
	full_add comp1747(.out(wire2599), .cout(wire2600), .inA(wire2300), .inB(wire2302), .cin(wire2304));
	full_add comp1748(.out(wire2601), .cout(wire2602), .inA(wire2305), .inB(wire2307), .cin(wire2309));
	full_add comp1749(.out(wire2603), .cout(wire2604), .inA(wire2306), .inB(wire2308), .cin(wire2310));
	full_add comp1750(.out(wire2605), .cout(wire2606), .inA(wire2311), .inB(wire2313), .cin(wire2315));
	full_add comp1751(.out(wire2607), .cout(wire2608), .inA(wire2312), .inB(wire2314), .cin(wire2316));
	full_add comp1752(.out(wire2609), .cout(wire2610), .inA(wire2317), .inB(wire2319), .cin(wire2321));
	full_add comp1753(.out(wire2611), .cout(wire2612), .inA(wire2318), .inB(wire2320), .cin(wire2322));
	full_add comp1754(.out(wire2613), .cout(wire2614), .inA(wire2323), .inB(wire2325), .cin(wire2327));
	full_add comp1755(.out(wire2615), .cout(wire2616), .inA(wire2324), .inB(wire2326), .cin(wire2328));
	full_add comp1756(.out(wire2617), .cout(wire2618), .inA(wire2329), .inB(wire2331), .cin(wire2333));
	full_add comp1757(.out(wire2619), .cout(wire2620), .inA(wire2330), .inB(wire2332), .cin(wire2334));
	full_add comp1758(.out(wire2621), .cout(wire2622), .inA(wire2335), .inB(wire2337), .cin(wire2339));
	full_add comp1759(.out(wire2623), .cout(wire2624), .inA(wire2336), .inB(wire2338), .cin(wire2340));
	full_add comp1760(.out(wire2625), .cout(wire2626), .inA(wire2341), .inB(wire2343), .cin(wire2345));
	full_add comp1761(.out(wire2627), .cout(wire2628), .inA(wire2342), .inB(wire2344), .cin(wire2346));
	full_add comp1762(.out(wire2629), .cout(wire2630), .inA(wire2347), .inB(wire2349), .cin(wire2351));
	full_add comp1763(.out(wire2631), .cout(wire2632), .inA(wire2348), .inB(wire2350), .cin(wire2352));
	full_add comp1764(.out(wire2633), .cout(wire2634), .inA(wire2353), .inB(wire2355), .cin(wire2357));
	full_add comp1765(.out(wire2635), .cout(wire2636), .inA(wire2354), .inB(wire2356), .cin(wire2358));
	full_add comp1766(.out(wire2637), .cout(wire2638), .inA(wire2359), .inB(wire2361), .cin(wire2363));
	full_add comp1767(.out(wire2639), .cout(wire2640), .inA(wire2360), .inB(wire2362), .cin(wire2364));
	full_add comp1768(.out(wire2641), .cout(wire2642), .inA(wire2365), .inB(wire2367), .cin(wire2369));
	full_add comp1769(.out(wire2643), .cout(wire2644), .inA(wire2366), .inB(wire2368), .cin(wire2370));
	full_add comp1770(.out(wire2645), .cout(wire2646), .inA(wire2371), .inB(wire2373), .cin(wire2375));
	full_add comp1771(.out(wire2647), .cout(wire2648), .inA(wire2372), .inB(wire2374), .cin(wire2376));
	full_add comp1772(.out(wire2649), .cout(wire2650), .inA(wire2377), .inB(wire2379), .cin(wire2381));
	full_add comp1773(.out(wire2651), .cout(wire2652), .inA(wire2378), .inB(wire2380), .cin(wire2382));
	full_add comp1774(.out(wire2653), .cout(wire2654), .inA(wire2383), .inB(wire2385), .cin(wire2387));
	full_add comp1775(.out(wire2655), .cout(wire2656), .inA(wire2384), .inB(wire2386), .cin(wire2388));
	full_add comp1776(.out(wire2657), .cout(wire2658), .inA(wire2389), .inB(wire2391), .cin(wire2393));
	full_add comp1777(.out(wire2659), .cout(wire2660), .inA(wire2390), .inB(wire2392), .cin(wire2394));
	full_add comp1778(.out(wire2661), .cout(wire2662), .inA(wire2395), .inB(wire2397), .cin(wire2399));
	full_add comp1779(.out(wire2663), .cout(wire2664), .inA(wire2396), .inB(wire2398), .cin(wire2400));
	full_add comp1780(.out(wire2665), .cout(wire2666), .inA(wire2401), .inB(wire2403), .cin(wire2405));
	full_add comp1781(.out(wire2667), .cout(wire2668), .inA(wire2402), .inB(wire2404), .cin(wire2406));
	full_add comp1782(.out(wire2669), .cout(wire2670), .inA(wire2407), .inB(wire2409), .cin(wire2411));
	full_add comp1783(.out(wire2671), .cout(wire2672), .inA(wire2408), .inB(wire2410), .cin(wire2412));
	full_add comp1784(.out(wire2673), .cout(wire2674), .inA(wire2413), .inB(wire2415), .cin(wire2417));
	full_add comp1785(.out(wire2675), .cout(wire2676), .inA(wire2414), .inB(wire2416), .cin(wire2418));
	full_add comp1786(.out(wire2677), .cout(wire2678), .inA(wire2419), .inB(wire2421), .cin(wire2423));
	full_add comp1787(.out(wire2679), .cout(wire2680), .inA(wire2420), .inB(wire2422), .cin(wire2424));
	full_add comp1788(.out(wire2681), .cout(wire2682), .inA(wire2425), .inB(wire2427), .cin(wire2429));
	full_add comp1789(.out(wire2683), .cout(wire2684), .inA(wire2426), .inB(wire2428), .cin(wire2430));
	full_add comp1790(.out(wire2685), .cout(wire2686), .inA(wire2431), .inB(wire2433), .cin(wire2435));
	full_add comp1791(.out(wire2687), .cout(wire2688), .inA(wire2432), .inB(wire2434), .cin(wire2436));
	full_add comp1792(.out(wire2689), .cout(wire2690), .inA(wire2437), .inB(wire2439), .cin(wire2441));
	full_add comp1793(.out(wire2691), .cout(wire2692), .inA(wire2438), .inB(wire2440), .cin(wire2442));
	full_add comp1794(.out(wire2693), .cout(wire2694), .inA(wire2443), .inB(wire2445), .cin(wire2447));
	full_add comp1795(.out(wire2695), .cout(wire2696), .inA(wire2444), .inB(wire2446), .cin(wire2448));
	full_add comp1796(.out(wire2697), .cout(wire2698), .inA(wire2449), .inB(wire2451), .cin(wire2453));
	full_add comp1797(.out(wire2699), .cout(wire2700), .inA(wire2450), .inB(wire2452), .cin(wire2454));
	full_add comp1798(.out(wire2701), .cout(wire2702), .inA(wire2455), .inB(wire2457), .cin(wire2459));
	full_add comp1799(.out(wire2703), .cout(wire2704), .inA(wire2456), .inB(wire2458), .cin(wire2460));
	full_add comp1800(.out(wire2705), .cout(wire2706), .inA(wire2461), .inB(wire2463), .cin(wire2465));
	full_add comp1801(.out(wire2707), .cout(wire2708), .inA(wire2462), .inB(wire2464), .cin(wire2466));
	full_add comp1802(.out(wire2709), .cout(wire2710), .inA(wire2467), .inB(wire2469), .cin(wire2471));
	full_add comp1803(.out(wire2711), .cout(wire2712), .inA(wire2468), .inB(wire2470), .cin(wire2472));
	full_add comp1804(.out(wire2713), .cout(wire2714), .inA(wire2473), .inB(wire2475), .cin(wire2477));
	full_add comp1805(.out(wire2715), .cout(wire2716), .inA(wire2474), .inB(wire2476), .cin(wire2478));
	full_add comp1806(.out(wire2717), .cout(wire2718), .inA(wire2479), .inB(wire2481), .cin(wire2483));
	full_add comp1807(.out(wire2719), .cout(wire2720), .inA(wire2480), .inB(wire2482), .cin(wire2484));
	full_add comp1808(.out(wire2721), .cout(wire2722), .inA(wire2485), .inB(wire2487), .cin(wire2489));
	full_add comp1809(.out(wire2723), .cout(wire2724), .inA(wire2486), .inB(wire2488), .cin(wire2490));
	full_add comp1810(.out(wire2725), .cout(wire2726), .inA(wire2491), .inB(wire2493), .cin(wire2495));
	full_add comp1811(.out(wire2727), .cout(wire2728), .inA(wire2492), .inB(wire2494), .cin(wire2496));
	full_add comp1812(.out(wire2729), .cout(wire2730), .inA(wire2497), .inB(wire2499), .cin(wire2501));
	full_add comp1813(.out(wire2731), .cout(wire2732), .inA(wire2498), .inB(wire2500), .cin(wire2502));
	full_add comp1814(.out(wire2733), .cout(wire2734), .inA(wire2503), .inB(wire2505), .cin(wire2507));
	full_add comp1815(.out(wire2735), .cout(wire2736), .inA(wire2504), .inB(wire2506), .cin(wire2508));
	full_add comp1816(.out(wire2737), .cout(wire2738), .inA(wire2509), .inB(wire2511), .cin(wire2513));
	full_add comp1817(.out(wire2739), .cout(wire2740), .inA(wire2510), .inB(wire2512), .cin(wire2514));
	full_add comp1818(.out(wire2741), .cout(wire2742), .inA(wire2515), .inB(wire2517), .cin(wire2519));
	full_add comp1819(.out(wire2743), .cout(wire2744), .inA(wire2516), .inB(wire2518), .cin(wire2520));
	full_add comp1820(.out(wire2745), .cout(wire2746), .inA(wire2521), .inB(wire2523), .cin(wire2525));
	full_add comp1821(.out(wire2747), .cout(wire2748), .inA(wire2522), .inB(wire2524), .cin(wire2526));
	full_add comp1822(.out(wire2749), .cout(wire2750), .inA(wire2527), .inB(wire2529), .cin(wire2531));
	full_add comp1823(.out(wire2751), .cout(wire2752), .inA(wire2528), .inB(wire2530), .cin(wire2532));
	full_add comp1824(.out(wire2753), .cout(wire2754), .inA(wire2533), .inB(wire2535), .cin(wire2537));
	full_add comp1825(.out(wire2755), .cout(wire2756), .inA(wire2534), .inB(wire2536), .cin(wire2538));
	full_add comp1826(.out(wire2757), .cout(wire2758), .inA(wire2539), .inB(wire2541), .cin(wire2543));
	full_add comp1827(.out(wire2759), .cout(wire2760), .inA(wire2540), .inB(wire2542), .cin(wire2544));
	full_add comp1828(.out(wire2761), .cout(wire2762), .inA(wire2545), .inB(wire2547), .cin(wire2549));
	full_add comp1829(.out(wire2763), .cout(wire2764), .inA(wire1146), .inB(wire2546), .cin(wire2548));
	full_add comp1830(.out(wire2765), .cout(wire2766), .inA(wire2550), .inB(wire2551), .cin(wire2553));
	full_add comp1831(.out(wire2767), .cout(wire2768), .inA(wire1085), .inB(wire1116), .cin(wire1147));
	full_add comp1832(.out(wire2769), .cout(wire2770), .inA(wire2552), .inB(wire2554), .cin(wire2555));
	full_add comp1833(.out(wire2771), .cout(wire2772), .inA(wire1024), .inB(wire1055), .cin(wire1086));
	full_add comp1834(.out(wire2773), .cout(wire2774), .inA(wire1117), .inB(wire1148), .cin(wire2556));
	full_add comp1835(.out(wire2775), .cout(wire2776), .inA(wire1056), .inB(wire1087), .cin(wire1118));
	half_add comp1836(.out(wire2777), .cout(wire2778), .inA(wire132), .inB(wire163));
	full_add comp1837(.out(wire2779), .cout(wire2780), .inA(wire195), .inB(wire226), .cin(wire257));
	full_add comp1838(.out(wire2781), .cout(wire2782), .inA(wire289), .inB(wire2558), .cin(wire2559));
	full_add comp1839(.out(wire2783), .cout(wire2784), .inA(wire2560), .inB(wire2562), .cin(wire2563));
	full_add comp1840(.out(wire2785), .cout(wire2786), .inA(wire2564), .inB(wire2566), .cin(wire2567));
	full_add comp1841(.out(wire2787), .cout(wire2788), .inA(wire2568), .inB(wire2570), .cin(wire2571));
	full_add comp1842(.out(wire2789), .cout(wire2790), .inA(wire2572), .inB(wire2574), .cin(wire2575));
	full_add comp1843(.out(wire2791), .cout(wire2792), .inA(wire2576), .inB(wire2578), .cin(wire2579));
	full_add comp1844(.out(wire2793), .cout(wire2794), .inA(wire2580), .inB(wire2582), .cin(wire2583));
	full_add comp1845(.out(wire2795), .cout(wire2796), .inA(wire2584), .inB(wire2586), .cin(wire2587));
	full_add comp1846(.out(wire2797), .cout(wire2798), .inA(wire2588), .inB(wire2590), .cin(wire2591));
	full_add comp1847(.out(wire2799), .cout(wire2800), .inA(wire2592), .inB(wire2594), .cin(wire2595));
	full_add comp1848(.out(wire2801), .cout(wire2802), .inA(wire2596), .inB(wire2598), .cin(wire2599));
	full_add comp1849(.out(wire2803), .cout(wire2804), .inA(wire2600), .inB(wire2602), .cin(wire2603));
	full_add comp1850(.out(wire2805), .cout(wire2806), .inA(wire2604), .inB(wire2606), .cin(wire2607));
	full_add comp1851(.out(wire2807), .cout(wire2808), .inA(wire2608), .inB(wire2610), .cin(wire2611));
	full_add comp1852(.out(wire2809), .cout(wire2810), .inA(wire2612), .inB(wire2614), .cin(wire2615));
	full_add comp1853(.out(wire2811), .cout(wire2812), .inA(wire2616), .inB(wire2618), .cin(wire2619));
	full_add comp1854(.out(wire2813), .cout(wire2814), .inA(wire2620), .inB(wire2622), .cin(wire2623));
	full_add comp1855(.out(wire2815), .cout(wire2816), .inA(wire2624), .inB(wire2626), .cin(wire2627));
	full_add comp1856(.out(wire2817), .cout(wire2818), .inA(wire2628), .inB(wire2630), .cin(wire2631));
	full_add comp1857(.out(wire2819), .cout(wire2820), .inA(wire2632), .inB(wire2634), .cin(wire2635));
	full_add comp1858(.out(wire2821), .cout(wire2822), .inA(wire2636), .inB(wire2638), .cin(wire2639));
	full_add comp1859(.out(wire2823), .cout(wire2824), .inA(wire2640), .inB(wire2642), .cin(wire2643));
	full_add comp1860(.out(wire2825), .cout(wire2826), .inA(wire2644), .inB(wire2646), .cin(wire2647));
	full_add comp1861(.out(wire2827), .cout(wire2828), .inA(wire2648), .inB(wire2650), .cin(wire2651));
	full_add comp1862(.out(wire2829), .cout(wire2830), .inA(wire2652), .inB(wire2654), .cin(wire2655));
	full_add comp1863(.out(wire2831), .cout(wire2832), .inA(wire2656), .inB(wire2658), .cin(wire2659));
	full_add comp1864(.out(wire2833), .cout(wire2834), .inA(wire2660), .inB(wire2662), .cin(wire2663));
	full_add comp1865(.out(wire2835), .cout(wire2836), .inA(wire2664), .inB(wire2666), .cin(wire2667));
	full_add comp1866(.out(wire2837), .cout(wire2838), .inA(wire2668), .inB(wire2670), .cin(wire2671));
	full_add comp1867(.out(wire2839), .cout(wire2840), .inA(wire2672), .inB(wire2674), .cin(wire2675));
	full_add comp1868(.out(wire2841), .cout(wire2842), .inA(wire2676), .inB(wire2678), .cin(wire2679));
	full_add comp1869(.out(wire2843), .cout(wire2844), .inA(wire2680), .inB(wire2682), .cin(wire2683));
	full_add comp1870(.out(wire2845), .cout(wire2846), .inA(wire2684), .inB(wire2686), .cin(wire2687));
	full_add comp1871(.out(wire2847), .cout(wire2848), .inA(wire2688), .inB(wire2690), .cin(wire2691));
	full_add comp1872(.out(wire2849), .cout(wire2850), .inA(wire2692), .inB(wire2694), .cin(wire2695));
	full_add comp1873(.out(wire2851), .cout(wire2852), .inA(wire2696), .inB(wire2698), .cin(wire2699));
	full_add comp1874(.out(wire2853), .cout(wire2854), .inA(wire2700), .inB(wire2702), .cin(wire2703));
	full_add comp1875(.out(wire2855), .cout(wire2856), .inA(wire2704), .inB(wire2706), .cin(wire2707));
	full_add comp1876(.out(wire2857), .cout(wire2858), .inA(wire2708), .inB(wire2710), .cin(wire2711));
	full_add comp1877(.out(wire2859), .cout(wire2860), .inA(wire2712), .inB(wire2714), .cin(wire2715));
	full_add comp1878(.out(wire2861), .cout(wire2862), .inA(wire2716), .inB(wire2718), .cin(wire2719));
	full_add comp1879(.out(wire2863), .cout(wire2864), .inA(wire2720), .inB(wire2722), .cin(wire2723));
	full_add comp1880(.out(wire2865), .cout(wire2866), .inA(wire2724), .inB(wire2726), .cin(wire2727));
	full_add comp1881(.out(wire2867), .cout(wire2868), .inA(wire2728), .inB(wire2730), .cin(wire2731));
	full_add comp1882(.out(wire2869), .cout(wire2870), .inA(wire2732), .inB(wire2734), .cin(wire2735));
	full_add comp1883(.out(wire2871), .cout(wire2872), .inA(wire2736), .inB(wire2738), .cin(wire2739));
	full_add comp1884(.out(wire2873), .cout(wire2874), .inA(wire2740), .inB(wire2742), .cin(wire2743));
	full_add comp1885(.out(wire2875), .cout(wire2876), .inA(wire2744), .inB(wire2746), .cin(wire2747));
	full_add comp1886(.out(wire2877), .cout(wire2878), .inA(wire2748), .inB(wire2750), .cin(wire2751));
	full_add comp1887(.out(wire2879), .cout(wire2880), .inA(wire2752), .inB(wire2754), .cin(wire2755));
	full_add comp1888(.out(wire2881), .cout(wire2882), .inA(wire2756), .inB(wire2758), .cin(wire2759));
	full_add comp1889(.out(wire2883), .cout(wire2884), .inA(wire2760), .inB(wire2762), .cin(wire2763));
	full_add comp1890(.out(wire2885), .cout(wire2886), .inA(wire2764), .inB(wire2766), .cin(wire2767));
	full_add comp1891(.out(wire2887), .cout(wire2888), .inA(wire2768), .inB(wire2770), .cin(wire2771));
	full_add comp1892(.out(wire2889), .cout(wire2890), .inA(wire1149), .inB(wire2772), .cin(wire2774));
	full_add comp1893(.out(wire2891), .cout(wire2892), .inA(wire1088), .inB(wire1119), .cin(wire1150));
	half_add comp1894(.out(wire2893), .cout(wire2894), .inA(wire131), .inB(wire162));
	full_add comp1895(.out(wire2895), .cout(wire2896), .inA(wire194), .inB(wire225), .cin(wire2777));
	full_add comp1896(.out(wire2897), .cout(wire2898), .inA(wire2557), .inB(wire2778), .cin(wire2779));
	full_add comp1897(.out(wire2899), .cout(wire2900), .inA(wire2561), .inB(wire2780), .cin(wire2781));
	full_add comp1898(.out(wire2901), .cout(wire2902), .inA(wire2565), .inB(wire2782), .cin(wire2783));
	full_add comp1899(.out(wire2903), .cout(wire2904), .inA(wire2569), .inB(wire2784), .cin(wire2785));
	full_add comp1900(.out(wire2905), .cout(wire2906), .inA(wire2573), .inB(wire2786), .cin(wire2787));
	full_add comp1901(.out(wire2907), .cout(wire2908), .inA(wire2577), .inB(wire2788), .cin(wire2789));
	full_add comp1902(.out(wire2909), .cout(wire2910), .inA(wire2581), .inB(wire2790), .cin(wire2791));
	full_add comp1903(.out(wire2911), .cout(wire2912), .inA(wire2585), .inB(wire2792), .cin(wire2793));
	full_add comp1904(.out(wire2913), .cout(wire2914), .inA(wire2589), .inB(wire2794), .cin(wire2795));
	full_add comp1905(.out(wire2915), .cout(wire2916), .inA(wire2593), .inB(wire2796), .cin(wire2797));
	full_add comp1906(.out(wire2917), .cout(wire2918), .inA(wire2597), .inB(wire2798), .cin(wire2799));
	full_add comp1907(.out(wire2919), .cout(wire2920), .inA(wire2601), .inB(wire2800), .cin(wire2801));
	full_add comp1908(.out(wire2921), .cout(wire2922), .inA(wire2605), .inB(wire2802), .cin(wire2803));
	full_add comp1909(.out(wire2923), .cout(wire2924), .inA(wire2609), .inB(wire2804), .cin(wire2805));
	full_add comp1910(.out(wire2925), .cout(wire2926), .inA(wire2613), .inB(wire2806), .cin(wire2807));
	full_add comp1911(.out(wire2927), .cout(wire2928), .inA(wire2617), .inB(wire2808), .cin(wire2809));
	full_add comp1912(.out(wire2929), .cout(wire2930), .inA(wire2621), .inB(wire2810), .cin(wire2811));
	full_add comp1913(.out(wire2931), .cout(wire2932), .inA(wire2625), .inB(wire2812), .cin(wire2813));
	full_add comp1914(.out(wire2933), .cout(wire2934), .inA(wire2629), .inB(wire2814), .cin(wire2815));
	full_add comp1915(.out(wire2935), .cout(wire2936), .inA(wire2633), .inB(wire2816), .cin(wire2817));
	full_add comp1916(.out(wire2937), .cout(wire2938), .inA(wire2637), .inB(wire2818), .cin(wire2819));
	full_add comp1917(.out(wire2939), .cout(wire2940), .inA(wire2641), .inB(wire2820), .cin(wire2821));
	full_add comp1918(.out(wire2941), .cout(wire2942), .inA(wire2645), .inB(wire2822), .cin(wire2823));
	full_add comp1919(.out(wire2943), .cout(wire2944), .inA(wire2649), .inB(wire2824), .cin(wire2825));
	full_add comp1920(.out(wire2945), .cout(wire2946), .inA(wire2653), .inB(wire2826), .cin(wire2827));
	full_add comp1921(.out(wire2947), .cout(wire2948), .inA(wire2657), .inB(wire2828), .cin(wire2829));
	full_add comp1922(.out(wire2949), .cout(wire2950), .inA(wire2661), .inB(wire2830), .cin(wire2831));
	full_add comp1923(.out(wire2951), .cout(wire2952), .inA(wire2665), .inB(wire2832), .cin(wire2833));
	full_add comp1924(.out(wire2953), .cout(wire2954), .inA(wire2669), .inB(wire2834), .cin(wire2835));
	full_add comp1925(.out(wire2955), .cout(wire2956), .inA(wire2673), .inB(wire2836), .cin(wire2837));
	full_add comp1926(.out(wire2957), .cout(wire2958), .inA(wire2677), .inB(wire2838), .cin(wire2839));
	full_add comp1927(.out(wire2959), .cout(wire2960), .inA(wire2681), .inB(wire2840), .cin(wire2841));
	full_add comp1928(.out(wire2961), .cout(wire2962), .inA(wire2685), .inB(wire2842), .cin(wire2843));
	full_add comp1929(.out(wire2963), .cout(wire2964), .inA(wire2689), .inB(wire2844), .cin(wire2845));
	full_add comp1930(.out(wire2965), .cout(wire2966), .inA(wire2693), .inB(wire2846), .cin(wire2847));
	full_add comp1931(.out(wire2967), .cout(wire2968), .inA(wire2697), .inB(wire2848), .cin(wire2849));
	full_add comp1932(.out(wire2969), .cout(wire2970), .inA(wire2701), .inB(wire2850), .cin(wire2851));
	full_add comp1933(.out(wire2971), .cout(wire2972), .inA(wire2705), .inB(wire2852), .cin(wire2853));
	full_add comp1934(.out(wire2973), .cout(wire2974), .inA(wire2709), .inB(wire2854), .cin(wire2855));
	full_add comp1935(.out(wire2975), .cout(wire2976), .inA(wire2713), .inB(wire2856), .cin(wire2857));
	full_add comp1936(.out(wire2977), .cout(wire2978), .inA(wire2717), .inB(wire2858), .cin(wire2859));
	full_add comp1937(.out(wire2979), .cout(wire2980), .inA(wire2721), .inB(wire2860), .cin(wire2861));
	full_add comp1938(.out(wire2981), .cout(wire2982), .inA(wire2725), .inB(wire2862), .cin(wire2863));
	full_add comp1939(.out(wire2983), .cout(wire2984), .inA(wire2729), .inB(wire2864), .cin(wire2865));
	full_add comp1940(.out(wire2985), .cout(wire2986), .inA(wire2733), .inB(wire2866), .cin(wire2867));
	full_add comp1941(.out(wire2987), .cout(wire2988), .inA(wire2737), .inB(wire2868), .cin(wire2869));
	full_add comp1942(.out(wire2989), .cout(wire2990), .inA(wire2741), .inB(wire2870), .cin(wire2871));
	full_add comp1943(.out(wire2991), .cout(wire2992), .inA(wire2745), .inB(wire2872), .cin(wire2873));
	full_add comp1944(.out(wire2993), .cout(wire2994), .inA(wire2749), .inB(wire2874), .cin(wire2875));
	full_add comp1945(.out(wire2995), .cout(wire2996), .inA(wire2753), .inB(wire2876), .cin(wire2877));
	full_add comp1946(.out(wire2997), .cout(wire2998), .inA(wire2757), .inB(wire2878), .cin(wire2879));
	full_add comp1947(.out(wire2999), .cout(wire3000), .inA(wire2761), .inB(wire2880), .cin(wire2881));
	full_add comp1948(.out(wire3001), .cout(wire3002), .inA(wire2765), .inB(wire2882), .cin(wire2883));
	full_add comp1949(.out(wire3003), .cout(wire3004), .inA(wire2769), .inB(wire2884), .cin(wire2885));
	full_add comp1950(.out(wire3005), .cout(wire3006), .inA(wire2773), .inB(wire2886), .cin(wire2887));
	full_add comp1951(.out(wire3007), .cout(wire3008), .inA(wire2775), .inB(wire2888), .cin(wire2889));
	full_add comp1952(.out(wire3009), .cout(wire3010), .inA(wire2776), .inB(wire2890), .cin(wire2891));
	full_add comp1953(.out(wire3011), .cout(wire3012), .inA(wire1120), .inB(wire1151), .cin(wire2892));
	wire [63:0] inA_comp1954;
	assign inA_comp1954[0] = wire129;
	assign inA_comp1954[1] = wire130;
	assign inA_comp1954[2] = wire193;
	assign inA_comp1954[3] = wire2894;
	assign inA_comp1954[4] = wire2896;
	assign inA_comp1954[5] = wire2898;
	assign inA_comp1954[6] = wire2900;
	assign inA_comp1954[7] = wire2902;
	assign inA_comp1954[8] = wire2904;
	assign inA_comp1954[9] = wire2906;
	assign inA_comp1954[10] = wire2908;
	assign inA_comp1954[11] = wire2910;
	assign inA_comp1954[12] = wire2912;
	assign inA_comp1954[13] = wire2914;
	assign inA_comp1954[14] = wire2916;
	assign inA_comp1954[15] = wire2918;
	assign inA_comp1954[16] = wire2920;
	assign inA_comp1954[17] = wire2922;
	assign inA_comp1954[18] = wire2924;
	assign inA_comp1954[19] = wire2926;
	assign inA_comp1954[20] = wire2928;
	assign inA_comp1954[21] = wire2930;
	assign inA_comp1954[22] = wire2932;
	assign inA_comp1954[23] = wire2934;
	assign inA_comp1954[24] = wire2936;
	assign inA_comp1954[25] = wire2938;
	assign inA_comp1954[26] = wire2940;
	assign inA_comp1954[27] = wire2942;
	assign inA_comp1954[28] = wire2944;
	assign inA_comp1954[29] = wire2946;
	assign inA_comp1954[30] = wire2948;
	assign inA_comp1954[31] = wire2950;
	assign inA_comp1954[32] = wire2952;
	assign inA_comp1954[33] = wire2954;
	assign inA_comp1954[34] = wire2956;
	assign inA_comp1954[35] = wire2958;
	assign inA_comp1954[36] = wire2960;
	assign inA_comp1954[37] = wire2962;
	assign inA_comp1954[38] = wire2964;
	assign inA_comp1954[39] = wire2966;
	assign inA_comp1954[40] = wire2968;
	assign inA_comp1954[41] = wire2970;
	assign inA_comp1954[42] = wire2972;
	assign inA_comp1954[43] = wire2974;
	assign inA_comp1954[44] = wire2976;
	assign inA_comp1954[45] = wire2978;
	assign inA_comp1954[46] = wire2980;
	assign inA_comp1954[47] = wire2982;
	assign inA_comp1954[48] = wire2984;
	assign inA_comp1954[49] = wire2986;
	assign inA_comp1954[50] = wire2988;
	assign inA_comp1954[51] = wire2990;
	assign inA_comp1954[52] = wire2992;
	assign inA_comp1954[53] = wire2994;
	assign inA_comp1954[54] = wire2996;
	assign inA_comp1954[55] = wire2998;
	assign inA_comp1954[56] = wire3000;
	assign inA_comp1954[57] = wire3002;
	assign inA_comp1954[58] = wire3004;
	assign inA_comp1954[59] = wire3006;
	assign inA_comp1954[60] = wire3008;
	assign inA_comp1954[61] = wire3010;
	assign inA_comp1954[62] = wire1152;
	assign inA_comp1954[63] = 1'b0;
	wire [63:0] inB_comp1954;
	assign inB_comp1954[0] = 1'b0;
	assign inB_comp1954[1] = wire161;
	assign inB_comp1954[2] = wire2893;
	assign inB_comp1954[3] = wire2895;
	assign inB_comp1954[4] = wire2897;
	assign inB_comp1954[5] = wire2899;
	assign inB_comp1954[6] = wire2901;
	assign inB_comp1954[7] = wire2903;
	assign inB_comp1954[8] = wire2905;
	assign inB_comp1954[9] = wire2907;
	assign inB_comp1954[10] = wire2909;
	assign inB_comp1954[11] = wire2911;
	assign inB_comp1954[12] = wire2913;
	assign inB_comp1954[13] = wire2915;
	assign inB_comp1954[14] = wire2917;
	assign inB_comp1954[15] = wire2919;
	assign inB_comp1954[16] = wire2921;
	assign inB_comp1954[17] = wire2923;
	assign inB_comp1954[18] = wire2925;
	assign inB_comp1954[19] = wire2927;
	assign inB_comp1954[20] = wire2929;
	assign inB_comp1954[21] = wire2931;
	assign inB_comp1954[22] = wire2933;
	assign inB_comp1954[23] = wire2935;
	assign inB_comp1954[24] = wire2937;
	assign inB_comp1954[25] = wire2939;
	assign inB_comp1954[26] = wire2941;
	assign inB_comp1954[27] = wire2943;
	assign inB_comp1954[28] = wire2945;
	assign inB_comp1954[29] = wire2947;
	assign inB_comp1954[30] = wire2949;
	assign inB_comp1954[31] = wire2951;
	assign inB_comp1954[32] = wire2953;
	assign inB_comp1954[33] = wire2955;
	assign inB_comp1954[34] = wire2957;
	assign inB_comp1954[35] = wire2959;
	assign inB_comp1954[36] = wire2961;
	assign inB_comp1954[37] = wire2963;
	assign inB_comp1954[38] = wire2965;
	assign inB_comp1954[39] = wire2967;
	assign inB_comp1954[40] = wire2969;
	assign inB_comp1954[41] = wire2971;
	assign inB_comp1954[42] = wire2973;
	assign inB_comp1954[43] = wire2975;
	assign inB_comp1954[44] = wire2977;
	assign inB_comp1954[45] = wire2979;
	assign inB_comp1954[46] = wire2981;
	assign inB_comp1954[47] = wire2983;
	assign inB_comp1954[48] = wire2985;
	assign inB_comp1954[49] = wire2987;
	assign inB_comp1954[50] = wire2989;
	assign inB_comp1954[51] = wire2991;
	assign inB_comp1954[52] = wire2993;
	assign inB_comp1954[53] = wire2995;
	assign inB_comp1954[54] = wire2997;
	assign inB_comp1954[55] = wire2999;
	assign inB_comp1954[56] = wire3001;
	assign inB_comp1954[57] = wire3003;
	assign inB_comp1954[58] = wire3005;
	assign inB_comp1954[59] = wire3007;
	assign inB_comp1954[60] = wire3009;
	assign inB_comp1954[61] = wire3011;
	assign inB_comp1954[62] = wire3012;
	assign inB_comp1954[63] = 1'b0;
	adder_64 comp1954(.out(out), .inA(inA_comp1954), .inB(inB_comp1954));

endmodule

